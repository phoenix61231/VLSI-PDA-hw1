
module GSIM_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  ADDHXL U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  ADDHXL U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  ADDHXL U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  ADDHXL U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  ADDHXL U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  ADDHXL U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  ADDHXL U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  ADDHXL U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  ADDHXL U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[31]), .B(A[31]), .Y(SUM[31]) );
endmodule


module GSIM_DW01_inc_1 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  ADDHXL U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  ADDHXL U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  ADDHXL U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  ADDHXL U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  ADDHXL U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  ADDHXL U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  ADDHXL U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  ADDHXL U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  ADDHXL U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  ADDHXL U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[31]), .B(A[31]), .Y(SUM[31]) );
endmodule


module GSIM_DW01_inc_2 ( A, SUM );
  input [63:0] A;
  output [63:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;

  NOR3BX1 U2 ( .AN(A[15]), .B(n12), .C(n72), .Y(n70) );
  NOR3BX1 U3 ( .AN(A[19]), .B(n11), .C(n68), .Y(n66) );
  NOR3BX1 U4 ( .AN(A[23]), .B(n10), .C(n64), .Y(n62) );
  NOR3BX1 U5 ( .AN(A[11]), .B(n13), .C(n76), .Y(n74) );
  NOR3BX1 U6 ( .AN(A[7]), .B(n14), .C(n19), .Y(n17) );
  NAND3X1 U7 ( .A(A[4]), .B(n26), .C(A[5]), .Y(n19) );
  NOR3BX1 U8 ( .AN(A[27]), .B(n9), .C(n60), .Y(n58) );
  NOR3BX1 U9 ( .AN(A[31]), .B(n8), .C(n56), .Y(n54) );
  NOR3BX1 U10 ( .AN(A[35]), .B(n7), .C(n52), .Y(n50) );
  NOR3BX1 U11 ( .AN(A[39]), .B(n6), .C(n46), .Y(n44) );
  NOR3BX1 U12 ( .AN(A[43]), .B(n5), .C(n42), .Y(n40) );
  NOR3BX1 U13 ( .AN(A[47]), .B(n4), .C(n38), .Y(n36) );
  NOR3BX1 U14 ( .AN(A[51]), .B(n3), .C(n34), .Y(n32) );
  NOR3BX1 U15 ( .AN(A[55]), .B(n2), .C(n30), .Y(n28) );
  NOR3BX1 U16 ( .AN(A[59]), .B(n1), .C(n24), .Y(n22) );
  NOR3BX1 U17 ( .AN(A[3]), .B(n15), .C(n48), .Y(n26) );
  XNOR2X1 U18 ( .A(A[61]), .B(n23), .Y(SUM[61]) );
  NOR2XL U19 ( .A(n24), .B(n1), .Y(n27) );
  NAND2XL U20 ( .A(A[56]), .B(n28), .Y(n29) );
  NOR2XL U21 ( .A(n30), .B(n2), .Y(n31) );
  NAND2XL U22 ( .A(A[52]), .B(n32), .Y(n33) );
  NOR2XL U23 ( .A(n34), .B(n3), .Y(n35) );
  NAND2XL U24 ( .A(A[48]), .B(n36), .Y(n37) );
  NOR2XL U25 ( .A(n38), .B(n4), .Y(n39) );
  NAND2XL U26 ( .A(A[44]), .B(n40), .Y(n41) );
  NOR2XL U27 ( .A(n42), .B(n5), .Y(n43) );
  NAND2XL U28 ( .A(A[40]), .B(n44), .Y(n45) );
  NOR2XL U29 ( .A(n46), .B(n6), .Y(n49) );
  NAND2XL U30 ( .A(A[36]), .B(n50), .Y(n51) );
  NOR2XL U31 ( .A(n52), .B(n7), .Y(n53) );
  NAND2XL U32 ( .A(A[32]), .B(n54), .Y(n55) );
  NOR2XL U33 ( .A(n56), .B(n8), .Y(n57) );
  NAND2XL U34 ( .A(A[28]), .B(n58), .Y(n59) );
  NOR2XL U35 ( .A(n60), .B(n9), .Y(n61) );
  NAND2XL U36 ( .A(A[24]), .B(n62), .Y(n63) );
  NOR2XL U37 ( .A(n64), .B(n10), .Y(n65) );
  NAND2XL U38 ( .A(A[20]), .B(n66), .Y(n67) );
  NOR2XL U39 ( .A(n68), .B(n11), .Y(n69) );
  NAND2XL U40 ( .A(A[16]), .B(n70), .Y(n71) );
  NOR2XL U41 ( .A(n72), .B(n12), .Y(n73) );
  NAND2XL U42 ( .A(A[12]), .B(n74), .Y(n75) );
  NOR2XL U43 ( .A(n76), .B(n13), .Y(n77) );
  NAND2XL U44 ( .A(A[8]), .B(n17), .Y(n16) );
  NOR2XL U45 ( .A(n19), .B(n14), .Y(n18) );
  NAND2XL U46 ( .A(A[4]), .B(n26), .Y(n25) );
  XOR2XL U47 ( .A(A[60]), .B(n22), .Y(SUM[60]) );
  NAND2XL U48 ( .A(A[60]), .B(n22), .Y(n23) );
  XNOR2XL U49 ( .A(A[62]), .B(n21), .Y(SUM[62]) );
  NOR2XL U50 ( .A(n48), .B(n15), .Y(n47) );
  CLKINVX1 U51 ( .A(A[58]), .Y(n1) );
  CLKINVX1 U52 ( .A(A[54]), .Y(n2) );
  CLKINVX1 U53 ( .A(A[50]), .Y(n3) );
  CLKINVX1 U54 ( .A(A[42]), .Y(n5) );
  CLKINVX1 U55 ( .A(A[38]), .Y(n6) );
  CLKINVX1 U56 ( .A(A[34]), .Y(n7) );
  CLKINVX1 U57 ( .A(A[30]), .Y(n8) );
  CLKINVX1 U58 ( .A(A[26]), .Y(n9) );
  CLKINVX1 U59 ( .A(A[46]), .Y(n4) );
  CLKINVX1 U60 ( .A(A[22]), .Y(n10) );
  CLKINVX1 U61 ( .A(A[18]), .Y(n11) );
  CLKINVX1 U62 ( .A(A[14]), .Y(n12) );
  CLKINVX1 U63 ( .A(A[10]), .Y(n13) );
  CLKINVX1 U64 ( .A(A[6]), .Y(n14) );
  CLKINVX1 U65 ( .A(A[2]), .Y(n15) );
  XNOR2X1 U66 ( .A(A[9]), .B(n16), .Y(SUM[9]) );
  XOR2X1 U67 ( .A(A[8]), .B(n17), .Y(SUM[8]) );
  XOR2X1 U68 ( .A(A[7]), .B(n18), .Y(SUM[7]) );
  XOR2X1 U69 ( .A(n14), .B(n19), .Y(SUM[6]) );
  XOR2X1 U70 ( .A(A[63]), .B(n20), .Y(SUM[63]) );
  NOR2BX1 U71 ( .AN(A[62]), .B(n21), .Y(n20) );
  NAND3X1 U72 ( .A(A[60]), .B(n22), .C(A[61]), .Y(n21) );
  XNOR2X1 U73 ( .A(A[5]), .B(n25), .Y(SUM[5]) );
  XOR2X1 U74 ( .A(A[59]), .B(n27), .Y(SUM[59]) );
  XOR2X1 U75 ( .A(n1), .B(n24), .Y(SUM[58]) );
  NAND3X1 U76 ( .A(A[56]), .B(n28), .C(A[57]), .Y(n24) );
  XNOR2X1 U77 ( .A(A[57]), .B(n29), .Y(SUM[57]) );
  XOR2X1 U78 ( .A(A[56]), .B(n28), .Y(SUM[56]) );
  XOR2X1 U79 ( .A(A[55]), .B(n31), .Y(SUM[55]) );
  XOR2X1 U80 ( .A(n2), .B(n30), .Y(SUM[54]) );
  NAND3X1 U81 ( .A(A[52]), .B(n32), .C(A[53]), .Y(n30) );
  XNOR2X1 U82 ( .A(A[53]), .B(n33), .Y(SUM[53]) );
  XOR2X1 U83 ( .A(A[52]), .B(n32), .Y(SUM[52]) );
  XOR2X1 U84 ( .A(A[51]), .B(n35), .Y(SUM[51]) );
  XOR2X1 U85 ( .A(n3), .B(n34), .Y(SUM[50]) );
  NAND3X1 U86 ( .A(A[48]), .B(n36), .C(A[49]), .Y(n34) );
  XOR2X1 U87 ( .A(A[4]), .B(n26), .Y(SUM[4]) );
  XNOR2X1 U88 ( .A(A[49]), .B(n37), .Y(SUM[49]) );
  XOR2X1 U89 ( .A(A[48]), .B(n36), .Y(SUM[48]) );
  XOR2X1 U90 ( .A(A[47]), .B(n39), .Y(SUM[47]) );
  XOR2X1 U91 ( .A(n4), .B(n38), .Y(SUM[46]) );
  NAND3X1 U92 ( .A(A[44]), .B(n40), .C(A[45]), .Y(n38) );
  XNOR2X1 U93 ( .A(A[45]), .B(n41), .Y(SUM[45]) );
  XOR2X1 U94 ( .A(A[44]), .B(n40), .Y(SUM[44]) );
  XOR2X1 U95 ( .A(A[43]), .B(n43), .Y(SUM[43]) );
  XOR2X1 U96 ( .A(n5), .B(n42), .Y(SUM[42]) );
  NAND3X1 U97 ( .A(A[40]), .B(n44), .C(A[41]), .Y(n42) );
  XNOR2X1 U98 ( .A(A[41]), .B(n45), .Y(SUM[41]) );
  XOR2X1 U99 ( .A(A[40]), .B(n44), .Y(SUM[40]) );
  XOR2X1 U100 ( .A(A[3]), .B(n47), .Y(SUM[3]) );
  XOR2X1 U101 ( .A(A[39]), .B(n49), .Y(SUM[39]) );
  XOR2X1 U102 ( .A(n6), .B(n46), .Y(SUM[38]) );
  NAND3X1 U103 ( .A(A[36]), .B(n50), .C(A[37]), .Y(n46) );
  XNOR2X1 U104 ( .A(A[37]), .B(n51), .Y(SUM[37]) );
  XOR2X1 U105 ( .A(A[36]), .B(n50), .Y(SUM[36]) );
  XOR2X1 U106 ( .A(A[35]), .B(n53), .Y(SUM[35]) );
  XOR2X1 U107 ( .A(n7), .B(n52), .Y(SUM[34]) );
  NAND3X1 U108 ( .A(A[32]), .B(n54), .C(A[33]), .Y(n52) );
  XNOR2X1 U109 ( .A(A[33]), .B(n55), .Y(SUM[33]) );
  XOR2X1 U110 ( .A(A[32]), .B(n54), .Y(SUM[32]) );
  XOR2X1 U111 ( .A(A[31]), .B(n57), .Y(SUM[31]) );
  XOR2X1 U112 ( .A(n8), .B(n56), .Y(SUM[30]) );
  NAND3X1 U113 ( .A(A[28]), .B(n58), .C(A[29]), .Y(n56) );
  XOR2X1 U114 ( .A(n15), .B(n48), .Y(SUM[2]) );
  XNOR2X1 U115 ( .A(A[29]), .B(n59), .Y(SUM[29]) );
  XOR2X1 U116 ( .A(A[28]), .B(n58), .Y(SUM[28]) );
  XOR2X1 U117 ( .A(A[27]), .B(n61), .Y(SUM[27]) );
  XOR2X1 U118 ( .A(n9), .B(n60), .Y(SUM[26]) );
  NAND3X1 U119 ( .A(A[24]), .B(n62), .C(A[25]), .Y(n60) );
  XNOR2X1 U120 ( .A(A[25]), .B(n63), .Y(SUM[25]) );
  XOR2X1 U121 ( .A(A[24]), .B(n62), .Y(SUM[24]) );
  XOR2X1 U122 ( .A(A[23]), .B(n65), .Y(SUM[23]) );
  XOR2X1 U123 ( .A(n10), .B(n64), .Y(SUM[22]) );
  NAND3X1 U124 ( .A(A[20]), .B(n66), .C(A[21]), .Y(n64) );
  XNOR2X1 U125 ( .A(A[21]), .B(n67), .Y(SUM[21]) );
  XOR2X1 U126 ( .A(A[20]), .B(n66), .Y(SUM[20]) );
  XOR2X1 U127 ( .A(A[19]), .B(n69), .Y(SUM[19]) );
  XOR2X1 U128 ( .A(n11), .B(n68), .Y(SUM[18]) );
  NAND3X1 U129 ( .A(A[16]), .B(n70), .C(A[17]), .Y(n68) );
  XNOR2X1 U130 ( .A(A[17]), .B(n71), .Y(SUM[17]) );
  XOR2X1 U131 ( .A(A[16]), .B(n70), .Y(SUM[16]) );
  XOR2X1 U132 ( .A(A[15]), .B(n73), .Y(SUM[15]) );
  XOR2X1 U133 ( .A(n12), .B(n72), .Y(SUM[14]) );
  NAND3X1 U134 ( .A(A[12]), .B(n74), .C(A[13]), .Y(n72) );
  XNOR2X1 U135 ( .A(A[13]), .B(n75), .Y(SUM[13]) );
  XOR2X1 U136 ( .A(A[12]), .B(n74), .Y(SUM[12]) );
  XOR2X1 U137 ( .A(A[11]), .B(n77), .Y(SUM[11]) );
  XOR2X1 U138 ( .A(n13), .B(n76), .Y(SUM[10]) );
  NAND3X1 U139 ( .A(A[8]), .B(n17), .C(A[9]), .Y(n76) );
  NAND2X1 U140 ( .A(A[1]), .B(A[0]), .Y(n48) );
endmodule


module GSIM_DW01_absval_0 ( A, ABSVAL );
  input [63:0] A;
  output [63:0] ABSVAL;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68;
  wire   [63:0] AMUX1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  GSIM_DW01_inc_2 NEG ( .A({n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
        n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
        n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
        n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
        n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68}), .SUM({
        AMUX1[63:2], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1}) );
  CLKINVX1 U1 ( .A(A[60]), .Y(n8) );
  CLKMX2X2 U2 ( .A(A[61]), .B(AMUX1[61]), .S0(n4), .Y(ABSVAL[61]) );
  CLKINVX1 U3 ( .A(A[62]), .Y(n6) );
  INVX3 U4 ( .A(n5), .Y(n4) );
  INVX3 U5 ( .A(n5), .Y(n3) );
  INVX3 U6 ( .A(n5), .Y(n2) );
  INVX3 U7 ( .A(n5), .Y(n1) );
  CLKINVX1 U8 ( .A(A[63]), .Y(n5) );
  CLKINVX1 U9 ( .A(A[58]), .Y(n10) );
  CLKINVX1 U10 ( .A(A[54]), .Y(n14) );
  CLKINVX1 U11 ( .A(A[57]), .Y(n11) );
  CLKINVX1 U12 ( .A(A[59]), .Y(n9) );
  CLKINVX1 U13 ( .A(A[55]), .Y(n13) );
  CLKINVX1 U14 ( .A(A[51]), .Y(n17) );
  CLKINVX1 U15 ( .A(A[47]), .Y(n21) );
  CLKINVX1 U16 ( .A(A[43]), .Y(n25) );
  CLKINVX1 U17 ( .A(A[56]), .Y(n12) );
  CLKINVX1 U18 ( .A(A[52]), .Y(n16) );
  CLKINVX1 U19 ( .A(A[48]), .Y(n20) );
  CLKINVX1 U20 ( .A(A[44]), .Y(n24) );
  CLKINVX1 U21 ( .A(A[50]), .Y(n18) );
  CLKINVX1 U22 ( .A(A[42]), .Y(n26) );
  CLKINVX1 U23 ( .A(A[38]), .Y(n30) );
  CLKINVX1 U24 ( .A(A[34]), .Y(n34) );
  CLKINVX1 U25 ( .A(A[30]), .Y(n38) );
  CLKINVX1 U26 ( .A(A[26]), .Y(n42) );
  CLKINVX1 U27 ( .A(A[61]), .Y(n7) );
  CLKINVX1 U28 ( .A(A[53]), .Y(n15) );
  CLKINVX1 U29 ( .A(A[49]), .Y(n19) );
  CLKINVX1 U30 ( .A(A[45]), .Y(n23) );
  CLKINVX1 U31 ( .A(A[41]), .Y(n27) );
  CLKINVX1 U32 ( .A(A[37]), .Y(n31) );
  CLKINVX1 U33 ( .A(A[33]), .Y(n35) );
  CLKINVX1 U34 ( .A(A[29]), .Y(n39) );
  CLKINVX1 U35 ( .A(A[39]), .Y(n29) );
  CLKINVX1 U36 ( .A(A[35]), .Y(n33) );
  CLKINVX1 U37 ( .A(A[31]), .Y(n37) );
  CLKINVX1 U38 ( .A(A[27]), .Y(n41) );
  CLKINVX1 U39 ( .A(A[23]), .Y(n45) );
  CLKINVX1 U40 ( .A(A[19]), .Y(n49) );
  CLKINVX1 U41 ( .A(A[15]), .Y(n53) );
  CLKINVX1 U42 ( .A(A[46]), .Y(n22) );
  CLKINVX1 U43 ( .A(A[40]), .Y(n28) );
  CLKINVX1 U44 ( .A(A[36]), .Y(n32) );
  CLKINVX1 U45 ( .A(A[32]), .Y(n36) );
  CLKINVX1 U46 ( .A(A[28]), .Y(n40) );
  CLKINVX1 U47 ( .A(A[24]), .Y(n44) );
  CLKINVX1 U48 ( .A(A[20]), .Y(n48) );
  CLKINVX1 U49 ( .A(A[16]), .Y(n52) );
  CLKINVX1 U50 ( .A(A[22]), .Y(n46) );
  CLKINVX1 U51 ( .A(A[18]), .Y(n50) );
  CLKINVX1 U52 ( .A(A[14]), .Y(n54) );
  CLKINVX1 U53 ( .A(A[10]), .Y(n58) );
  CLKINVX1 U54 ( .A(A[6]), .Y(n62) );
  CLKINVX1 U55 ( .A(A[2]), .Y(n66) );
  CLKINVX1 U56 ( .A(A[25]), .Y(n43) );
  CLKINVX1 U57 ( .A(A[21]), .Y(n47) );
  CLKINVX1 U58 ( .A(A[17]), .Y(n51) );
  CLKINVX1 U59 ( .A(A[13]), .Y(n55) );
  CLKINVX1 U60 ( .A(A[9]), .Y(n59) );
  CLKINVX1 U61 ( .A(A[5]), .Y(n63) );
  CLKINVX1 U62 ( .A(A[11]), .Y(n57) );
  CLKINVX1 U63 ( .A(A[7]), .Y(n61) );
  CLKINVX1 U64 ( .A(A[3]), .Y(n65) );
  CLKINVX1 U65 ( .A(A[12]), .Y(n56) );
  CLKINVX1 U66 ( .A(A[8]), .Y(n60) );
  CLKINVX1 U67 ( .A(A[4]), .Y(n64) );
  CLKINVX1 U68 ( .A(A[0]), .Y(n68) );
  CLKINVX1 U69 ( .A(A[1]), .Y(n67) );
  CLKMX2X2 U70 ( .A(A[9]), .B(AMUX1[9]), .S0(n3), .Y(ABSVAL[9]) );
  CLKMX2X2 U71 ( .A(A[8]), .B(AMUX1[8]), .S0(n4), .Y(ABSVAL[8]) );
  CLKMX2X2 U72 ( .A(A[7]), .B(AMUX1[7]), .S0(n4), .Y(ABSVAL[7]) );
  CLKMX2X2 U73 ( .A(A[6]), .B(AMUX1[6]), .S0(n4), .Y(ABSVAL[6]) );
  AND2X1 U74 ( .A(AMUX1[63]), .B(n4), .Y(ABSVAL[63]) );
  CLKMX2X2 U75 ( .A(A[62]), .B(AMUX1[62]), .S0(n4), .Y(ABSVAL[62]) );
  CLKMX2X2 U76 ( .A(A[60]), .B(AMUX1[60]), .S0(n4), .Y(ABSVAL[60]) );
  CLKMX2X2 U77 ( .A(A[5]), .B(AMUX1[5]), .S0(n4), .Y(ABSVAL[5]) );
  CLKMX2X2 U78 ( .A(A[59]), .B(AMUX1[59]), .S0(n4), .Y(ABSVAL[59]) );
  CLKMX2X2 U79 ( .A(A[58]), .B(AMUX1[58]), .S0(n4), .Y(ABSVAL[58]) );
  CLKMX2X2 U80 ( .A(A[57]), .B(AMUX1[57]), .S0(n4), .Y(ABSVAL[57]) );
  CLKMX2X2 U81 ( .A(A[56]), .B(AMUX1[56]), .S0(n3), .Y(ABSVAL[56]) );
  CLKMX2X2 U82 ( .A(A[55]), .B(AMUX1[55]), .S0(n3), .Y(ABSVAL[55]) );
  CLKMX2X2 U83 ( .A(A[54]), .B(AMUX1[54]), .S0(n3), .Y(ABSVAL[54]) );
  CLKMX2X2 U84 ( .A(A[53]), .B(AMUX1[53]), .S0(n3), .Y(ABSVAL[53]) );
  CLKMX2X2 U85 ( .A(A[52]), .B(AMUX1[52]), .S0(n3), .Y(ABSVAL[52]) );
  CLKMX2X2 U86 ( .A(A[51]), .B(AMUX1[51]), .S0(n3), .Y(ABSVAL[51]) );
  CLKMX2X2 U87 ( .A(A[50]), .B(AMUX1[50]), .S0(n3), .Y(ABSVAL[50]) );
  CLKMX2X2 U88 ( .A(A[4]), .B(AMUX1[4]), .S0(n3), .Y(ABSVAL[4]) );
  CLKMX2X2 U89 ( .A(A[49]), .B(AMUX1[49]), .S0(n3), .Y(ABSVAL[49]) );
  CLKMX2X2 U90 ( .A(A[48]), .B(AMUX1[48]), .S0(n3), .Y(ABSVAL[48]) );
  CLKMX2X2 U91 ( .A(A[47]), .B(AMUX1[47]), .S0(n3), .Y(ABSVAL[47]) );
  CLKMX2X2 U92 ( .A(A[46]), .B(AMUX1[46]), .S0(n3), .Y(ABSVAL[46]) );
  CLKMX2X2 U93 ( .A(A[45]), .B(AMUX1[45]), .S0(n3), .Y(ABSVAL[45]) );
  CLKMX2X2 U94 ( .A(A[44]), .B(AMUX1[44]), .S0(n2), .Y(ABSVAL[44]) );
  CLKMX2X2 U95 ( .A(A[43]), .B(AMUX1[43]), .S0(n2), .Y(ABSVAL[43]) );
  CLKMX2X2 U96 ( .A(A[42]), .B(AMUX1[42]), .S0(n2), .Y(ABSVAL[42]) );
  CLKMX2X2 U97 ( .A(A[41]), .B(AMUX1[41]), .S0(n2), .Y(ABSVAL[41]) );
  CLKMX2X2 U98 ( .A(A[40]), .B(AMUX1[40]), .S0(n2), .Y(ABSVAL[40]) );
  CLKMX2X2 U99 ( .A(A[3]), .B(AMUX1[3]), .S0(n2), .Y(ABSVAL[3]) );
  CLKMX2X2 U100 ( .A(A[39]), .B(AMUX1[39]), .S0(n2), .Y(ABSVAL[39]) );
  CLKMX2X2 U101 ( .A(A[38]), .B(AMUX1[38]), .S0(n2), .Y(ABSVAL[38]) );
  CLKMX2X2 U102 ( .A(A[37]), .B(AMUX1[37]), .S0(n2), .Y(ABSVAL[37]) );
  CLKMX2X2 U103 ( .A(A[36]), .B(AMUX1[36]), .S0(n2), .Y(ABSVAL[36]) );
  CLKMX2X2 U104 ( .A(A[35]), .B(AMUX1[35]), .S0(n2), .Y(ABSVAL[35]) );
  CLKMX2X2 U105 ( .A(A[34]), .B(AMUX1[34]), .S0(n2), .Y(ABSVAL[34]) );
  CLKMX2X2 U106 ( .A(A[33]), .B(AMUX1[33]), .S0(n1), .Y(ABSVAL[33]) );
  CLKMX2X2 U107 ( .A(A[32]), .B(AMUX1[32]), .S0(n1), .Y(ABSVAL[32]) );
  CLKMX2X2 U108 ( .A(A[31]), .B(AMUX1[31]), .S0(n1), .Y(ABSVAL[31]) );
  CLKMX2X2 U109 ( .A(A[30]), .B(AMUX1[30]), .S0(n1), .Y(ABSVAL[30]) );
  CLKMX2X2 U110 ( .A(A[2]), .B(AMUX1[2]), .S0(n1), .Y(ABSVAL[2]) );
  CLKMX2X2 U111 ( .A(A[29]), .B(AMUX1[29]), .S0(n1), .Y(ABSVAL[29]) );
  CLKMX2X2 U112 ( .A(A[28]), .B(AMUX1[28]), .S0(n1), .Y(ABSVAL[28]) );
  CLKMX2X2 U113 ( .A(A[27]), .B(AMUX1[27]), .S0(n1), .Y(ABSVAL[27]) );
  CLKMX2X2 U114 ( .A(A[26]), .B(AMUX1[26]), .S0(n1), .Y(ABSVAL[26]) );
  CLKMX2X2 U115 ( .A(A[25]), .B(AMUX1[25]), .S0(n1), .Y(ABSVAL[25]) );
  CLKMX2X2 U116 ( .A(A[24]), .B(AMUX1[24]), .S0(n1), .Y(ABSVAL[24]) );
  CLKMX2X2 U117 ( .A(A[23]), .B(AMUX1[23]), .S0(n1), .Y(ABSVAL[23]) );
  CLKMX2X2 U118 ( .A(A[22]), .B(AMUX1[22]), .S0(n1), .Y(ABSVAL[22]) );
  CLKMX2X2 U119 ( .A(A[21]), .B(AMUX1[21]), .S0(n1), .Y(ABSVAL[21]) );
  CLKMX2X2 U120 ( .A(A[20]), .B(AMUX1[20]), .S0(n1), .Y(ABSVAL[20]) );
  CLKMX2X2 U121 ( .A(A[19]), .B(AMUX1[19]), .S0(n1), .Y(ABSVAL[19]) );
  CLKMX2X2 U122 ( .A(A[18]), .B(AMUX1[18]), .S0(n1), .Y(ABSVAL[18]) );
  CLKMX2X2 U123 ( .A(A[17]), .B(AMUX1[17]), .S0(n2), .Y(ABSVAL[17]) );
  CLKMX2X2 U124 ( .A(A[16]), .B(AMUX1[16]), .S0(n2), .Y(ABSVAL[16]) );
  CLKMX2X2 U125 ( .A(A[15]), .B(AMUX1[15]), .S0(n2), .Y(ABSVAL[15]) );
  CLKMX2X2 U126 ( .A(A[14]), .B(AMUX1[14]), .S0(n2), .Y(ABSVAL[14]) );
  CLKMX2X2 U127 ( .A(A[13]), .B(AMUX1[13]), .S0(n3), .Y(ABSVAL[13]) );
  CLKMX2X2 U128 ( .A(A[12]), .B(AMUX1[12]), .S0(n3), .Y(ABSVAL[12]) );
  CLKMX2X2 U129 ( .A(A[11]), .B(AMUX1[11]), .S0(n3), .Y(ABSVAL[11]) );
  CLKMX2X2 U130 ( .A(A[10]), .B(AMUX1[10]), .S0(n2), .Y(ABSVAL[10]) );
endmodule


module GSIM_DW_inc_0 ( carry_in, a, carry_out, sum );
  input [63:0] a;
  output [63:0] sum;
  input carry_in;
  output carry_out;
  wire   \sum[63] , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63;
  assign sum[62] = \sum[63] ;
  assign sum[61] = \sum[63] ;
  assign sum[63] = \sum[63] ;

  ADDHXL U7 ( .A(a[59]), .B(n5), .CO(n4), .S(sum[59]) );
  ADDHXL U9 ( .A(a[57]), .B(n7), .CO(n6), .S(sum[57]) );
  ADDHXL U12 ( .A(a[54]), .B(n10), .CO(n9), .S(sum[54]) );
  ADDHXL U15 ( .A(a[51]), .B(n13), .CO(n12), .S(sum[51]) );
  ADDHXL U19 ( .A(a[47]), .B(n17), .CO(n16), .S(sum[47]) );
  ADDHXL U22 ( .A(a[44]), .B(n20), .CO(n19), .S(sum[44]) );
  ADDHXL U25 ( .A(a[41]), .B(n23), .CO(n22), .S(sum[41]) );
  ADDHXL U30 ( .A(a[36]), .B(n28), .CO(n27), .S(sum[36]) );
  ADDHXL U33 ( .A(a[33]), .B(n31), .CO(n30), .S(sum[33]) );
  ADDHXL U35 ( .A(a[31]), .B(n33), .CO(n32), .S(sum[31]) );
  ADDHXL U41 ( .A(a[25]), .B(n39), .CO(n38), .S(sum[25]) );
  ADDHXL U44 ( .A(a[22]), .B(n42), .CO(n41), .S(sum[22]) );
  ADDHXL U46 ( .A(a[20]), .B(n44), .CO(n43), .S(sum[20]) );
  ADDHXL U50 ( .A(a[16]), .B(n48), .CO(n47), .S(sum[16]) );
  ADDHXL U52 ( .A(a[14]), .B(n50), .CO(n49), .S(sum[14]) );
  ADDHXL U54 ( .A(a[12]), .B(n52), .CO(n51), .S(sum[12]) );
  ADDHXL U56 ( .A(a[10]), .B(n54), .CO(n53), .S(sum[10]) );
  ADDHXL U60 ( .A(a[6]), .B(n58), .CO(n57), .S(sum[6]) );
  ADDHXL U62 ( .A(a[4]), .B(n60), .CO(n59), .S(sum[4]) );
  ADDHXL U66 ( .A(carry_in), .B(a[0]), .CO(n63), .S(sum[0]) );
  ADDHX2 U70 ( .A(a[2]), .B(n62), .CO(n61), .S(sum[2]) );
  ADDHX2 U71 ( .A(a[1]), .B(n63), .CO(n62), .S(sum[1]) );
  ADDHXL U72 ( .A(a[11]), .B(n53), .CO(n52), .S(sum[11]) );
  ADDHXL U73 ( .A(a[13]), .B(n51), .CO(n50), .S(sum[13]) );
  ADDHXL U74 ( .A(a[15]), .B(n49), .CO(n48), .S(sum[15]) );
  ADDHXL U75 ( .A(a[17]), .B(n47), .CO(n46), .S(sum[17]) );
  ADDHXL U76 ( .A(a[19]), .B(n45), .CO(n44), .S(sum[19]) );
  ADDHXL U77 ( .A(a[23]), .B(n41), .CO(n40), .S(sum[23]) );
  ADDHXL U78 ( .A(a[21]), .B(n43), .CO(n42), .S(sum[21]) );
  ADDHXL U79 ( .A(a[5]), .B(n59), .CO(n58), .S(sum[5]) );
  ADDHXL U80 ( .A(a[9]), .B(n55), .CO(n54), .S(sum[9]) );
  ADDHXL U81 ( .A(a[3]), .B(n61), .CO(n60), .S(sum[3]) );
  ADDHXL U82 ( .A(a[7]), .B(n57), .CO(n56), .S(sum[7]) );
  ADDHXL U83 ( .A(a[26]), .B(n38), .CO(n37), .S(sum[26]) );
  ADDHXL U84 ( .A(a[29]), .B(n35), .CO(n34), .S(sum[29]) );
  ADDHXL U85 ( .A(a[32]), .B(n32), .CO(n31), .S(sum[32]) );
  ADDHXL U86 ( .A(a[34]), .B(n30), .CO(n29), .S(sum[34]) );
  ADDHXL U87 ( .A(a[37]), .B(n27), .CO(n26), .S(sum[37]) );
  ADDHXL U88 ( .A(a[39]), .B(n25), .CO(n24), .S(sum[39]) );
  ADDHXL U89 ( .A(a[42]), .B(n22), .CO(n21), .S(sum[42]) );
  ADDHXL U90 ( .A(a[45]), .B(n19), .CO(n18), .S(sum[45]) );
  ADDHXL U91 ( .A(a[48]), .B(n16), .CO(n15), .S(sum[48]) );
  ADDHXL U92 ( .A(a[50]), .B(n14), .CO(n13), .S(sum[50]) );
  ADDHXL U93 ( .A(a[52]), .B(n12), .CO(n11), .S(sum[52]) );
  ADDHXL U94 ( .A(a[53]), .B(n11), .CO(n10), .S(sum[53]) );
  ADDHXL U95 ( .A(a[55]), .B(n9), .CO(n8), .S(sum[55]) );
  ADDHXL U96 ( .A(a[56]), .B(n8), .CO(n7), .S(sum[56]) );
  ADDHXL U97 ( .A(a[58]), .B(n6), .CO(n5), .S(sum[58]) );
  ADDHXL U98 ( .A(a[35]), .B(n29), .CO(n28), .S(sum[35]) );
  ADDHXL U99 ( .A(a[24]), .B(n40), .CO(n39), .S(sum[24]) );
  ADDHXL U100 ( .A(a[43]), .B(n21), .CO(n20), .S(sum[43]) );
  ADDHXL U101 ( .A(a[27]), .B(n37), .CO(n36), .S(sum[27]) );
  ADDHXL U102 ( .A(a[46]), .B(n18), .CO(n17), .S(sum[46]) );
  ADDHXL U103 ( .A(a[30]), .B(n34), .CO(n33), .S(sum[30]) );
  ADDHXL U104 ( .A(a[40]), .B(n24), .CO(n23), .S(sum[40]) );
  NOR2BX1 U105 ( .AN(a[60]), .B(n4), .Y(\sum[63] ) );
  XOR2XL U106 ( .A(n4), .B(a[60]), .Y(sum[60]) );
  ADDHXL U107 ( .A(a[28]), .B(n36), .CO(n35), .S(sum[28]) );
  ADDHXL U108 ( .A(a[38]), .B(n26), .CO(n25), .S(sum[38]) );
  ADDHXL U109 ( .A(a[8]), .B(n56), .CO(n55), .S(sum[8]) );
  ADDHXL U110 ( .A(a[18]), .B(n46), .CO(n45), .S(sum[18]) );
  ADDHXL U111 ( .A(a[49]), .B(n15), .CO(n14), .S(sum[49]) );
endmodule


module GSIM_DW_div_tc_0 ( a, b, quotient, remainder, divide_by_0 );
  input [63:0] a;
  input [5:0] b;
  output [63:0] quotient;
  output [5:0] remainder;
  output divide_by_0;
  wire   \u_div/QInv[63] , \u_div/QInv[59] , \u_div/QInv[58] ,
         \u_div/QInv[57] , \u_div/QInv[56] , \u_div/QInv[55] ,
         \u_div/QInv[54] , \u_div/QInv[53] , \u_div/QInv[52] ,
         \u_div/QInv[51] , \u_div/QInv[50] , \u_div/QInv[49] ,
         \u_div/QInv[48] , \u_div/QInv[47] , \u_div/QInv[46] ,
         \u_div/QInv[45] , \u_div/QInv[44] , \u_div/QInv[43] ,
         \u_div/QInv[42] , \u_div/QInv[41] , \u_div/QInv[40] ,
         \u_div/QInv[39] , \u_div/QInv[38] , \u_div/QInv[37] ,
         \u_div/QInv[36] , \u_div/QInv[35] , \u_div/QInv[34] ,
         \u_div/QInv[33] , \u_div/QInv[32] , \u_div/QInv[31] ,
         \u_div/QInv[30] , \u_div/QInv[29] , \u_div/QInv[28] ,
         \u_div/QInv[27] , \u_div/QInv[26] , \u_div/QInv[25] ,
         \u_div/QInv[24] , \u_div/QInv[23] , \u_div/QInv[22] ,
         \u_div/QInv[21] , \u_div/QInv[20] , \u_div/QInv[19] ,
         \u_div/QInv[18] , \u_div/QInv[17] , \u_div/QInv[16] ,
         \u_div/QInv[15] , \u_div/QInv[14] , \u_div/QInv[13] ,
         \u_div/QInv[12] , \u_div/QInv[11] , \u_div/QInv[10] , \u_div/QInv[9] ,
         \u_div/QInv[8] , \u_div/QInv[7] , \u_div/QInv[6] , \u_div/QInv[5] ,
         \u_div/QInv[4] , \u_div/QInv[3] , \u_div/QInv[2] , \u_div/QInv[1] ,
         \u_div/QInv[0] , \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] ,
         \u_div/SumTmp[1][3] , \u_div/SumTmp[1][4] , \u_div/SumTmp[2][1] ,
         \u_div/SumTmp[2][2] , \u_div/SumTmp[2][3] , \u_div/SumTmp[2][4] ,
         \u_div/SumTmp[3][1] , \u_div/SumTmp[3][2] , \u_div/SumTmp[3][3] ,
         \u_div/SumTmp[3][4] , \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] ,
         \u_div/SumTmp[4][3] , \u_div/SumTmp[4][4] , \u_div/SumTmp[5][1] ,
         \u_div/SumTmp[5][2] , \u_div/SumTmp[5][3] , \u_div/SumTmp[5][4] ,
         \u_div/SumTmp[6][1] , \u_div/SumTmp[6][2] , \u_div/SumTmp[6][3] ,
         \u_div/SumTmp[6][4] , \u_div/SumTmp[7][1] , \u_div/SumTmp[7][2] ,
         \u_div/SumTmp[7][3] , \u_div/SumTmp[7][4] , \u_div/SumTmp[8][1] ,
         \u_div/SumTmp[8][2] , \u_div/SumTmp[8][3] , \u_div/SumTmp[8][4] ,
         \u_div/SumTmp[9][1] , \u_div/SumTmp[9][2] , \u_div/SumTmp[9][3] ,
         \u_div/SumTmp[9][4] , \u_div/SumTmp[10][1] , \u_div/SumTmp[10][2] ,
         \u_div/SumTmp[10][3] , \u_div/SumTmp[10][4] , \u_div/SumTmp[11][1] ,
         \u_div/SumTmp[11][2] , \u_div/SumTmp[11][3] , \u_div/SumTmp[11][4] ,
         \u_div/SumTmp[12][1] , \u_div/SumTmp[12][2] , \u_div/SumTmp[12][3] ,
         \u_div/SumTmp[12][4] , \u_div/SumTmp[13][1] , \u_div/SumTmp[13][2] ,
         \u_div/SumTmp[13][3] , \u_div/SumTmp[13][4] , \u_div/SumTmp[14][1] ,
         \u_div/SumTmp[14][2] , \u_div/SumTmp[14][3] , \u_div/SumTmp[14][4] ,
         \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] , \u_div/SumTmp[15][3] ,
         \u_div/SumTmp[15][4] , \u_div/SumTmp[16][1] , \u_div/SumTmp[16][2] ,
         \u_div/SumTmp[16][3] , \u_div/SumTmp[16][4] , \u_div/SumTmp[17][1] ,
         \u_div/SumTmp[17][2] , \u_div/SumTmp[17][3] , \u_div/SumTmp[17][4] ,
         \u_div/SumTmp[18][1] , \u_div/SumTmp[18][2] , \u_div/SumTmp[18][3] ,
         \u_div/SumTmp[18][4] , \u_div/SumTmp[19][1] , \u_div/SumTmp[19][2] ,
         \u_div/SumTmp[19][3] , \u_div/SumTmp[19][4] , \u_div/SumTmp[20][1] ,
         \u_div/SumTmp[20][2] , \u_div/SumTmp[20][3] , \u_div/SumTmp[20][4] ,
         \u_div/SumTmp[21][1] , \u_div/SumTmp[21][2] , \u_div/SumTmp[21][3] ,
         \u_div/SumTmp[21][4] , \u_div/SumTmp[22][1] , \u_div/SumTmp[22][2] ,
         \u_div/SumTmp[22][3] , \u_div/SumTmp[22][4] , \u_div/SumTmp[23][1] ,
         \u_div/SumTmp[23][2] , \u_div/SumTmp[23][3] , \u_div/SumTmp[23][4] ,
         \u_div/SumTmp[24][1] , \u_div/SumTmp[24][2] , \u_div/SumTmp[24][3] ,
         \u_div/SumTmp[24][4] , \u_div/SumTmp[25][1] , \u_div/SumTmp[25][2] ,
         \u_div/SumTmp[25][3] , \u_div/SumTmp[25][4] , \u_div/SumTmp[26][1] ,
         \u_div/SumTmp[26][2] , \u_div/SumTmp[26][3] , \u_div/SumTmp[26][4] ,
         \u_div/SumTmp[27][1] , \u_div/SumTmp[27][2] , \u_div/SumTmp[27][3] ,
         \u_div/SumTmp[27][4] , \u_div/SumTmp[28][1] , \u_div/SumTmp[28][2] ,
         \u_div/SumTmp[28][3] , \u_div/SumTmp[28][4] , \u_div/SumTmp[29][1] ,
         \u_div/SumTmp[29][2] , \u_div/SumTmp[29][3] , \u_div/SumTmp[29][4] ,
         \u_div/SumTmp[30][1] , \u_div/SumTmp[30][2] , \u_div/SumTmp[30][3] ,
         \u_div/SumTmp[30][4] , \u_div/SumTmp[31][1] , \u_div/SumTmp[31][2] ,
         \u_div/SumTmp[31][3] , \u_div/SumTmp[31][4] , \u_div/SumTmp[32][1] ,
         \u_div/SumTmp[32][2] , \u_div/SumTmp[32][3] , \u_div/SumTmp[32][4] ,
         \u_div/SumTmp[33][1] , \u_div/SumTmp[33][2] , \u_div/SumTmp[33][3] ,
         \u_div/SumTmp[33][4] , \u_div/SumTmp[34][1] , \u_div/SumTmp[34][2] ,
         \u_div/SumTmp[34][3] , \u_div/SumTmp[34][4] , \u_div/SumTmp[35][1] ,
         \u_div/SumTmp[35][2] , \u_div/SumTmp[35][3] , \u_div/SumTmp[35][4] ,
         \u_div/SumTmp[36][1] , \u_div/SumTmp[36][2] , \u_div/SumTmp[36][3] ,
         \u_div/SumTmp[36][4] , \u_div/SumTmp[37][1] , \u_div/SumTmp[37][2] ,
         \u_div/SumTmp[37][3] , \u_div/SumTmp[37][4] , \u_div/SumTmp[38][1] ,
         \u_div/SumTmp[38][2] , \u_div/SumTmp[38][3] , \u_div/SumTmp[38][4] ,
         \u_div/SumTmp[39][1] , \u_div/SumTmp[39][2] , \u_div/SumTmp[39][3] ,
         \u_div/SumTmp[39][4] , \u_div/SumTmp[40][1] , \u_div/SumTmp[40][2] ,
         \u_div/SumTmp[40][3] , \u_div/SumTmp[40][4] , \u_div/SumTmp[41][1] ,
         \u_div/SumTmp[41][2] , \u_div/SumTmp[41][3] , \u_div/SumTmp[41][4] ,
         \u_div/SumTmp[42][1] , \u_div/SumTmp[42][2] , \u_div/SumTmp[42][3] ,
         \u_div/SumTmp[42][4] , \u_div/SumTmp[43][1] , \u_div/SumTmp[43][2] ,
         \u_div/SumTmp[43][3] , \u_div/SumTmp[43][4] , \u_div/SumTmp[44][1] ,
         \u_div/SumTmp[44][2] , \u_div/SumTmp[44][3] , \u_div/SumTmp[44][4] ,
         \u_div/SumTmp[45][1] , \u_div/SumTmp[45][2] , \u_div/SumTmp[45][3] ,
         \u_div/SumTmp[45][4] , \u_div/SumTmp[46][1] , \u_div/SumTmp[46][2] ,
         \u_div/SumTmp[46][3] , \u_div/SumTmp[46][4] , \u_div/SumTmp[47][1] ,
         \u_div/SumTmp[47][2] , \u_div/SumTmp[47][3] , \u_div/SumTmp[47][4] ,
         \u_div/SumTmp[48][1] , \u_div/SumTmp[48][2] , \u_div/SumTmp[48][3] ,
         \u_div/SumTmp[48][4] , \u_div/SumTmp[49][1] , \u_div/SumTmp[49][2] ,
         \u_div/SumTmp[49][3] , \u_div/SumTmp[49][4] , \u_div/SumTmp[50][1] ,
         \u_div/SumTmp[50][2] , \u_div/SumTmp[50][3] , \u_div/SumTmp[50][4] ,
         \u_div/SumTmp[51][1] , \u_div/SumTmp[51][2] , \u_div/SumTmp[51][3] ,
         \u_div/SumTmp[51][4] , \u_div/SumTmp[52][1] , \u_div/SumTmp[52][2] ,
         \u_div/SumTmp[52][3] , \u_div/SumTmp[52][4] , \u_div/SumTmp[53][1] ,
         \u_div/SumTmp[53][2] , \u_div/SumTmp[53][3] , \u_div/SumTmp[53][4] ,
         \u_div/SumTmp[54][1] , \u_div/SumTmp[54][2] , \u_div/SumTmp[54][3] ,
         \u_div/SumTmp[54][4] , \u_div/SumTmp[55][1] , \u_div/SumTmp[55][2] ,
         \u_div/SumTmp[55][3] , \u_div/SumTmp[55][4] , \u_div/SumTmp[56][1] ,
         \u_div/SumTmp[56][2] , \u_div/SumTmp[56][3] , \u_div/SumTmp[56][4] ,
         \u_div/SumTmp[57][1] , \u_div/SumTmp[57][2] , \u_div/SumTmp[57][3] ,
         \u_div/SumTmp[57][4] , \u_div/SumTmp[58][1] , \u_div/SumTmp[58][2] ,
         \u_div/SumTmp[58][3] , \u_div/SumTmp[58][4] , \u_div/SumTmp[59][3] ,
         \u_div/SumTmp[59][4] , \u_div/CryTmp[0][6] , \u_div/CryTmp[1][6] ,
         \u_div/CryTmp[2][6] , \u_div/CryTmp[3][6] , \u_div/CryTmp[4][6] ,
         \u_div/CryTmp[5][6] , \u_div/CryTmp[6][6] , \u_div/CryTmp[7][6] ,
         \u_div/CryTmp[8][6] , \u_div/CryTmp[9][6] , \u_div/CryTmp[10][6] ,
         \u_div/CryTmp[11][6] , \u_div/CryTmp[12][6] , \u_div/CryTmp[13][6] ,
         \u_div/CryTmp[14][6] , \u_div/CryTmp[15][6] , \u_div/CryTmp[16][6] ,
         \u_div/CryTmp[17][6] , \u_div/CryTmp[18][6] , \u_div/CryTmp[19][6] ,
         \u_div/CryTmp[20][6] , \u_div/CryTmp[21][6] , \u_div/CryTmp[22][6] ,
         \u_div/CryTmp[23][6] , \u_div/CryTmp[24][6] , \u_div/CryTmp[25][6] ,
         \u_div/CryTmp[26][6] , \u_div/CryTmp[27][6] , \u_div/CryTmp[28][6] ,
         \u_div/CryTmp[29][6] , \u_div/CryTmp[30][6] , \u_div/CryTmp[31][6] ,
         \u_div/CryTmp[32][6] , \u_div/CryTmp[33][6] , \u_div/CryTmp[34][6] ,
         \u_div/CryTmp[35][6] , \u_div/CryTmp[36][6] , \u_div/CryTmp[37][6] ,
         \u_div/CryTmp[38][6] , \u_div/CryTmp[39][6] , \u_div/CryTmp[40][6] ,
         \u_div/CryTmp[41][6] , \u_div/CryTmp[42][6] , \u_div/CryTmp[43][6] ,
         \u_div/CryTmp[44][6] , \u_div/CryTmp[45][6] , \u_div/CryTmp[46][6] ,
         \u_div/CryTmp[47][6] , \u_div/CryTmp[48][6] , \u_div/CryTmp[49][6] ,
         \u_div/CryTmp[50][6] , \u_div/CryTmp[51][6] , \u_div/CryTmp[52][6] ,
         \u_div/CryTmp[53][6] , \u_div/CryTmp[54][6] , \u_div/CryTmp[55][6] ,
         \u_div/CryTmp[56][6] , \u_div/CryTmp[57][6] , \u_div/CryTmp[58][6] ,
         \u_div/CryTmp[59][6] , \u_div/PartRem[1][3] , \u_div/PartRem[1][4] ,
         \u_div/PartRem[1][5] , \u_div/PartRem[2][2] , \u_div/PartRem[2][3] ,
         \u_div/PartRem[2][4] , \u_div/PartRem[2][5] , \u_div/PartRem[3][0] ,
         \u_div/PartRem[3][2] , \u_div/PartRem[3][3] , \u_div/PartRem[3][4] ,
         \u_div/PartRem[3][5] , \u_div/PartRem[4][0] , \u_div/PartRem[4][2] ,
         \u_div/PartRem[4][3] , \u_div/PartRem[4][4] , \u_div/PartRem[4][5] ,
         \u_div/PartRem[5][0] , \u_div/PartRem[5][2] , \u_div/PartRem[5][3] ,
         \u_div/PartRem[5][4] , \u_div/PartRem[5][5] , \u_div/PartRem[6][0] ,
         \u_div/PartRem[6][2] , \u_div/PartRem[6][3] , \u_div/PartRem[6][4] ,
         \u_div/PartRem[6][5] , \u_div/PartRem[7][0] , \u_div/PartRem[7][2] ,
         \u_div/PartRem[7][3] , \u_div/PartRem[7][4] , \u_div/PartRem[7][5] ,
         \u_div/PartRem[8][0] , \u_div/PartRem[8][2] , \u_div/PartRem[8][3] ,
         \u_div/PartRem[8][4] , \u_div/PartRem[8][5] , \u_div/PartRem[9][0] ,
         \u_div/PartRem[9][2] , \u_div/PartRem[9][3] , \u_div/PartRem[9][4] ,
         \u_div/PartRem[9][5] , \u_div/PartRem[10][0] , \u_div/PartRem[10][2] ,
         \u_div/PartRem[10][3] , \u_div/PartRem[10][4] ,
         \u_div/PartRem[10][5] , \u_div/PartRem[11][0] ,
         \u_div/PartRem[11][2] , \u_div/PartRem[11][3] ,
         \u_div/PartRem[11][4] , \u_div/PartRem[11][5] ,
         \u_div/PartRem[12][0] , \u_div/PartRem[12][2] ,
         \u_div/PartRem[12][3] , \u_div/PartRem[12][4] ,
         \u_div/PartRem[12][5] , \u_div/PartRem[13][0] ,
         \u_div/PartRem[13][2] , \u_div/PartRem[13][3] ,
         \u_div/PartRem[13][4] , \u_div/PartRem[13][5] ,
         \u_div/PartRem[14][0] , \u_div/PartRem[14][2] ,
         \u_div/PartRem[14][3] , \u_div/PartRem[14][4] ,
         \u_div/PartRem[14][5] , \u_div/PartRem[15][0] ,
         \u_div/PartRem[15][2] , \u_div/PartRem[15][3] ,
         \u_div/PartRem[15][4] , \u_div/PartRem[15][5] ,
         \u_div/PartRem[16][0] , \u_div/PartRem[16][2] ,
         \u_div/PartRem[16][3] , \u_div/PartRem[16][4] ,
         \u_div/PartRem[16][5] , \u_div/PartRem[17][0] ,
         \u_div/PartRem[17][2] , \u_div/PartRem[17][3] ,
         \u_div/PartRem[17][4] , \u_div/PartRem[17][5] ,
         \u_div/PartRem[18][0] , \u_div/PartRem[18][2] ,
         \u_div/PartRem[18][3] , \u_div/PartRem[18][4] ,
         \u_div/PartRem[18][5] , \u_div/PartRem[19][0] ,
         \u_div/PartRem[19][2] , \u_div/PartRem[19][3] ,
         \u_div/PartRem[19][4] , \u_div/PartRem[19][5] ,
         \u_div/PartRem[20][0] , \u_div/PartRem[20][2] ,
         \u_div/PartRem[20][3] , \u_div/PartRem[20][4] ,
         \u_div/PartRem[20][5] , \u_div/PartRem[21][0] ,
         \u_div/PartRem[21][2] , \u_div/PartRem[21][3] ,
         \u_div/PartRem[21][4] , \u_div/PartRem[21][5] ,
         \u_div/PartRem[22][0] , \u_div/PartRem[22][2] ,
         \u_div/PartRem[22][3] , \u_div/PartRem[22][4] ,
         \u_div/PartRem[22][5] , \u_div/PartRem[23][0] ,
         \u_div/PartRem[23][2] , \u_div/PartRem[23][3] ,
         \u_div/PartRem[23][4] , \u_div/PartRem[23][5] ,
         \u_div/PartRem[24][0] , \u_div/PartRem[24][2] ,
         \u_div/PartRem[24][3] , \u_div/PartRem[24][4] ,
         \u_div/PartRem[24][5] , \u_div/PartRem[25][0] ,
         \u_div/PartRem[25][2] , \u_div/PartRem[25][3] ,
         \u_div/PartRem[25][4] , \u_div/PartRem[25][5] ,
         \u_div/PartRem[26][0] , \u_div/PartRem[26][2] ,
         \u_div/PartRem[26][3] , \u_div/PartRem[26][4] ,
         \u_div/PartRem[26][5] , \u_div/PartRem[27][0] ,
         \u_div/PartRem[27][2] , \u_div/PartRem[27][3] ,
         \u_div/PartRem[27][4] , \u_div/PartRem[27][5] ,
         \u_div/PartRem[28][0] , \u_div/PartRem[28][2] ,
         \u_div/PartRem[28][3] , \u_div/PartRem[28][4] ,
         \u_div/PartRem[28][5] , \u_div/PartRem[29][0] ,
         \u_div/PartRem[29][2] , \u_div/PartRem[29][3] ,
         \u_div/PartRem[29][4] , \u_div/PartRem[29][5] ,
         \u_div/PartRem[30][0] , \u_div/PartRem[30][2] ,
         \u_div/PartRem[30][3] , \u_div/PartRem[30][4] ,
         \u_div/PartRem[30][5] , \u_div/PartRem[31][0] ,
         \u_div/PartRem[31][2] , \u_div/PartRem[31][3] ,
         \u_div/PartRem[31][4] , \u_div/PartRem[31][5] ,
         \u_div/PartRem[32][0] , \u_div/PartRem[32][2] ,
         \u_div/PartRem[32][3] , \u_div/PartRem[32][4] ,
         \u_div/PartRem[32][5] , \u_div/PartRem[33][0] ,
         \u_div/PartRem[33][2] , \u_div/PartRem[33][3] ,
         \u_div/PartRem[33][4] , \u_div/PartRem[33][5] ,
         \u_div/PartRem[34][0] , \u_div/PartRem[34][2] ,
         \u_div/PartRem[34][3] , \u_div/PartRem[34][4] ,
         \u_div/PartRem[34][5] , \u_div/PartRem[35][0] ,
         \u_div/PartRem[35][2] , \u_div/PartRem[35][3] ,
         \u_div/PartRem[35][4] , \u_div/PartRem[35][5] ,
         \u_div/PartRem[36][0] , \u_div/PartRem[36][2] ,
         \u_div/PartRem[36][3] , \u_div/PartRem[36][4] ,
         \u_div/PartRem[36][5] , \u_div/PartRem[37][0] ,
         \u_div/PartRem[37][2] , \u_div/PartRem[37][3] ,
         \u_div/PartRem[37][4] , \u_div/PartRem[37][5] ,
         \u_div/PartRem[38][0] , \u_div/PartRem[38][2] ,
         \u_div/PartRem[38][3] , \u_div/PartRem[38][4] ,
         \u_div/PartRem[38][5] , \u_div/PartRem[39][0] ,
         \u_div/PartRem[39][2] , \u_div/PartRem[39][3] ,
         \u_div/PartRem[39][4] , \u_div/PartRem[39][5] ,
         \u_div/PartRem[40][0] , \u_div/PartRem[40][2] ,
         \u_div/PartRem[40][3] , \u_div/PartRem[40][4] ,
         \u_div/PartRem[40][5] , \u_div/PartRem[41][0] ,
         \u_div/PartRem[41][2] , \u_div/PartRem[41][3] ,
         \u_div/PartRem[41][4] , \u_div/PartRem[41][5] ,
         \u_div/PartRem[42][0] , \u_div/PartRem[42][2] ,
         \u_div/PartRem[42][3] , \u_div/PartRem[42][4] ,
         \u_div/PartRem[42][5] , \u_div/PartRem[43][0] ,
         \u_div/PartRem[43][2] , \u_div/PartRem[43][3] ,
         \u_div/PartRem[43][4] , \u_div/PartRem[43][5] ,
         \u_div/PartRem[44][0] , \u_div/PartRem[44][2] ,
         \u_div/PartRem[44][3] , \u_div/PartRem[44][4] ,
         \u_div/PartRem[44][5] , \u_div/PartRem[45][0] ,
         \u_div/PartRem[45][2] , \u_div/PartRem[45][3] ,
         \u_div/PartRem[45][4] , \u_div/PartRem[45][5] ,
         \u_div/PartRem[46][0] , \u_div/PartRem[46][2] ,
         \u_div/PartRem[46][3] , \u_div/PartRem[46][4] ,
         \u_div/PartRem[46][5] , \u_div/PartRem[47][0] ,
         \u_div/PartRem[47][2] , \u_div/PartRem[47][3] ,
         \u_div/PartRem[47][4] , \u_div/PartRem[47][5] ,
         \u_div/PartRem[48][0] , \u_div/PartRem[48][2] ,
         \u_div/PartRem[48][3] , \u_div/PartRem[48][4] ,
         \u_div/PartRem[48][5] , \u_div/PartRem[49][0] ,
         \u_div/PartRem[49][2] , \u_div/PartRem[49][3] ,
         \u_div/PartRem[49][4] , \u_div/PartRem[49][5] ,
         \u_div/PartRem[50][0] , \u_div/PartRem[50][2] ,
         \u_div/PartRem[50][3] , \u_div/PartRem[50][4] ,
         \u_div/PartRem[50][5] , \u_div/PartRem[51][0] ,
         \u_div/PartRem[51][2] , \u_div/PartRem[51][3] ,
         \u_div/PartRem[51][4] , \u_div/PartRem[51][5] ,
         \u_div/PartRem[52][0] , \u_div/PartRem[52][2] ,
         \u_div/PartRem[52][3] , \u_div/PartRem[52][4] ,
         \u_div/PartRem[52][5] , \u_div/PartRem[53][0] ,
         \u_div/PartRem[53][2] , \u_div/PartRem[53][3] ,
         \u_div/PartRem[53][4] , \u_div/PartRem[53][5] ,
         \u_div/PartRem[54][0] , \u_div/PartRem[54][2] ,
         \u_div/PartRem[54][3] , \u_div/PartRem[54][4] ,
         \u_div/PartRem[54][5] , \u_div/PartRem[55][0] ,
         \u_div/PartRem[55][2] , \u_div/PartRem[55][3] ,
         \u_div/PartRem[55][4] , \u_div/PartRem[55][5] ,
         \u_div/PartRem[56][0] , \u_div/PartRem[56][2] ,
         \u_div/PartRem[56][3] , \u_div/PartRem[56][4] ,
         \u_div/PartRem[56][5] , \u_div/PartRem[57][0] ,
         \u_div/PartRem[57][2] , \u_div/PartRem[57][3] ,
         \u_div/PartRem[57][4] , \u_div/PartRem[57][5] ,
         \u_div/PartRem[58][0] , \u_div/PartRem[58][2] ,
         \u_div/PartRem[58][3] , \u_div/PartRem[58][4] ,
         \u_div/PartRem[58][5] , \u_div/PartRem[59][0] ,
         \u_div/PartRem[59][2] , \u_div/PartRem[59][3] ,
         \u_div/PartRem[59][4] , \u_div/PartRem[59][5] ,
         \u_div/PartRem[60][0] , \u_div/PartRem[61][0] ,
         \u_div/PartRem[62][0] , \u_div/PartRem[63][0] ,
         \u_div/PartRem[64][0] , \u_div/u_add_PartRem_2_1/n3 ,
         \u_div/u_add_PartRem_2_1/n2 , \u_div/u_add_PartRem_2_2/n3 ,
         \u_div/u_add_PartRem_2_2/n2 , \u_div/u_add_PartRem_2_3/n3 ,
         \u_div/u_add_PartRem_2_3/n2 , \u_div/u_add_PartRem_2_4/n3 ,
         \u_div/u_add_PartRem_2_4/n2 , \u_div/u_add_PartRem_2_5/n3 ,
         \u_div/u_add_PartRem_2_5/n2 , \u_div/u_add_PartRem_2_6/n3 ,
         \u_div/u_add_PartRem_2_6/n2 , \u_div/u_add_PartRem_2_7/n3 ,
         \u_div/u_add_PartRem_2_7/n2 , \u_div/u_add_PartRem_2_8/n3 ,
         \u_div/u_add_PartRem_2_8/n2 , \u_div/u_add_PartRem_2_9/n3 ,
         \u_div/u_add_PartRem_2_9/n2 , \u_div/u_add_PartRem_2_10/n3 ,
         \u_div/u_add_PartRem_2_10/n2 , \u_div/u_add_PartRem_2_11/n3 ,
         \u_div/u_add_PartRem_2_11/n2 , \u_div/u_add_PartRem_2_12/n3 ,
         \u_div/u_add_PartRem_2_12/n2 , \u_div/u_add_PartRem_2_13/n3 ,
         \u_div/u_add_PartRem_2_13/n2 , \u_div/u_add_PartRem_2_14/n3 ,
         \u_div/u_add_PartRem_2_14/n2 , \u_div/u_add_PartRem_2_15/n3 ,
         \u_div/u_add_PartRem_2_15/n2 , \u_div/u_add_PartRem_2_16/n3 ,
         \u_div/u_add_PartRem_2_16/n2 , \u_div/u_add_PartRem_2_17/n3 ,
         \u_div/u_add_PartRem_2_17/n2 , \u_div/u_add_PartRem_2_18/n3 ,
         \u_div/u_add_PartRem_2_18/n2 , \u_div/u_add_PartRem_2_19/n3 ,
         \u_div/u_add_PartRem_2_19/n2 , \u_div/u_add_PartRem_2_20/n3 ,
         \u_div/u_add_PartRem_2_20/n2 , \u_div/u_add_PartRem_2_21/n3 ,
         \u_div/u_add_PartRem_2_21/n2 , \u_div/u_add_PartRem_2_22/n3 ,
         \u_div/u_add_PartRem_2_22/n2 , \u_div/u_add_PartRem_2_23/n3 ,
         \u_div/u_add_PartRem_2_23/n2 , \u_div/u_add_PartRem_2_24/n3 ,
         \u_div/u_add_PartRem_2_24/n2 , \u_div/u_add_PartRem_2_25/n3 ,
         \u_div/u_add_PartRem_2_25/n2 , \u_div/u_add_PartRem_2_26/n3 ,
         \u_div/u_add_PartRem_2_26/n2 , \u_div/u_add_PartRem_2_27/n3 ,
         \u_div/u_add_PartRem_2_27/n2 , \u_div/u_add_PartRem_2_28/n3 ,
         \u_div/u_add_PartRem_2_28/n2 , \u_div/u_add_PartRem_2_29/n3 ,
         \u_div/u_add_PartRem_2_29/n2 , \u_div/u_add_PartRem_2_30/n3 ,
         \u_div/u_add_PartRem_2_30/n2 , \u_div/u_add_PartRem_2_31/n3 ,
         \u_div/u_add_PartRem_2_31/n2 , \u_div/u_add_PartRem_2_32/n3 ,
         \u_div/u_add_PartRem_2_32/n2 , \u_div/u_add_PartRem_2_33/n3 ,
         \u_div/u_add_PartRem_2_33/n2 , \u_div/u_add_PartRem_2_34/n3 ,
         \u_div/u_add_PartRem_2_34/n2 , \u_div/u_add_PartRem_2_35/n3 ,
         \u_div/u_add_PartRem_2_35/n2 , \u_div/u_add_PartRem_2_36/n3 ,
         \u_div/u_add_PartRem_2_36/n2 , \u_div/u_add_PartRem_2_37/n3 ,
         \u_div/u_add_PartRem_2_37/n2 , \u_div/u_add_PartRem_2_38/n3 ,
         \u_div/u_add_PartRem_2_38/n2 , \u_div/u_add_PartRem_2_39/n3 ,
         \u_div/u_add_PartRem_2_39/n2 , \u_div/u_add_PartRem_2_40/n3 ,
         \u_div/u_add_PartRem_2_40/n2 , \u_div/u_add_PartRem_2_41/n3 ,
         \u_div/u_add_PartRem_2_41/n2 , \u_div/u_add_PartRem_2_42/n3 ,
         \u_div/u_add_PartRem_2_42/n2 , \u_div/u_add_PartRem_2_43/n3 ,
         \u_div/u_add_PartRem_2_43/n2 , \u_div/u_add_PartRem_2_44/n3 ,
         \u_div/u_add_PartRem_2_44/n2 , \u_div/u_add_PartRem_2_45/n3 ,
         \u_div/u_add_PartRem_2_45/n2 , \u_div/u_add_PartRem_2_46/n3 ,
         \u_div/u_add_PartRem_2_46/n2 , \u_div/u_add_PartRem_2_47/n3 ,
         \u_div/u_add_PartRem_2_47/n2 , \u_div/u_add_PartRem_2_48/n3 ,
         \u_div/u_add_PartRem_2_48/n2 , \u_div/u_add_PartRem_2_49/n3 ,
         \u_div/u_add_PartRem_2_49/n2 , \u_div/u_add_PartRem_2_50/n3 ,
         \u_div/u_add_PartRem_2_50/n2 , \u_div/u_add_PartRem_2_51/n3 ,
         \u_div/u_add_PartRem_2_51/n2 , \u_div/u_add_PartRem_2_52/n3 ,
         \u_div/u_add_PartRem_2_52/n2 , \u_div/u_add_PartRem_2_53/n3 ,
         \u_div/u_add_PartRem_2_53/n2 , \u_div/u_add_PartRem_2_54/n3 ,
         \u_div/u_add_PartRem_2_54/n2 , \u_div/u_add_PartRem_2_55/n3 ,
         \u_div/u_add_PartRem_2_55/n2 , \u_div/u_add_PartRem_2_56/n3 ,
         \u_div/u_add_PartRem_2_56/n2 , \u_div/u_add_PartRem_2_57/n3 ,
         \u_div/u_add_PartRem_2_57/n2 , \u_div/u_add_PartRem_2_58/n3 ,
         \u_div/u_add_PartRem_2_58/n2 , n1, n2, n3, n4, n5, n6, n7, n8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign \u_div/QInv[63]  = a[63];

  GSIM_DW01_absval_0 \u_div/u_absval_AAbs  ( .A({n3, a[62:0]}), .ABSVAL({
        \u_div/PartRem[64][0] , \u_div/PartRem[63][0] , \u_div/PartRem[62][0] , 
        \u_div/PartRem[61][0] , \u_div/PartRem[60][0] , \u_div/PartRem[59][0] , 
        \u_div/PartRem[58][0] , \u_div/PartRem[57][0] , \u_div/PartRem[56][0] , 
        \u_div/PartRem[55][0] , \u_div/PartRem[54][0] , \u_div/PartRem[53][0] , 
        \u_div/PartRem[52][0] , \u_div/PartRem[51][0] , \u_div/PartRem[50][0] , 
        \u_div/PartRem[49][0] , \u_div/PartRem[48][0] , \u_div/PartRem[47][0] , 
        \u_div/PartRem[46][0] , \u_div/PartRem[45][0] , \u_div/PartRem[44][0] , 
        \u_div/PartRem[43][0] , \u_div/PartRem[42][0] , \u_div/PartRem[41][0] , 
        \u_div/PartRem[40][0] , \u_div/PartRem[39][0] , \u_div/PartRem[38][0] , 
        \u_div/PartRem[37][0] , \u_div/PartRem[36][0] , \u_div/PartRem[35][0] , 
        \u_div/PartRem[34][0] , \u_div/PartRem[33][0] , \u_div/PartRem[32][0] , 
        \u_div/PartRem[31][0] , \u_div/PartRem[30][0] , \u_div/PartRem[29][0] , 
        \u_div/PartRem[28][0] , \u_div/PartRem[27][0] , \u_div/PartRem[26][0] , 
        \u_div/PartRem[25][0] , \u_div/PartRem[24][0] , \u_div/PartRem[23][0] , 
        \u_div/PartRem[22][0] , \u_div/PartRem[21][0] , \u_div/PartRem[20][0] , 
        \u_div/PartRem[19][0] , \u_div/PartRem[18][0] , \u_div/PartRem[17][0] , 
        \u_div/PartRem[16][0] , \u_div/PartRem[15][0] , \u_div/PartRem[14][0] , 
        \u_div/PartRem[13][0] , \u_div/PartRem[12][0] , \u_div/PartRem[11][0] , 
        \u_div/PartRem[10][0] , \u_div/PartRem[9][0] , \u_div/PartRem[8][0] , 
        \u_div/PartRem[7][0] , \u_div/PartRem[6][0] , \u_div/PartRem[5][0] , 
        \u_div/PartRem[4][0] , \u_div/PartRem[3][0] , SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1}) );
  GSIM_DW_inc_0 \u_div/u_inc_QInc  ( .carry_in(n4), .a({n3, n3, n3, 
        \u_div/QInv[63] , \u_div/QInv[59] , \u_div/QInv[58] , \u_div/QInv[57] , 
        \u_div/QInv[56] , \u_div/QInv[55] , \u_div/QInv[54] , \u_div/QInv[53] , 
        \u_div/QInv[52] , \u_div/QInv[51] , \u_div/QInv[50] , \u_div/QInv[49] , 
        \u_div/QInv[48] , \u_div/QInv[47] , \u_div/QInv[46] , \u_div/QInv[45] , 
        \u_div/QInv[44] , \u_div/QInv[43] , \u_div/QInv[42] , \u_div/QInv[41] , 
        \u_div/QInv[40] , \u_div/QInv[39] , \u_div/QInv[38] , \u_div/QInv[37] , 
        \u_div/QInv[36] , \u_div/QInv[35] , \u_div/QInv[34] , \u_div/QInv[33] , 
        \u_div/QInv[32] , \u_div/QInv[31] , \u_div/QInv[30] , \u_div/QInv[29] , 
        \u_div/QInv[28] , \u_div/QInv[27] , \u_div/QInv[26] , \u_div/QInv[25] , 
        \u_div/QInv[24] , \u_div/QInv[23] , \u_div/QInv[22] , \u_div/QInv[21] , 
        \u_div/QInv[20] , \u_div/QInv[19] , \u_div/QInv[18] , \u_div/QInv[17] , 
        \u_div/QInv[16] , \u_div/QInv[15] , \u_div/QInv[14] , \u_div/QInv[13] , 
        \u_div/QInv[12] , \u_div/QInv[11] , \u_div/QInv[10] , \u_div/QInv[9] , 
        \u_div/QInv[8] , \u_div/QInv[7] , \u_div/QInv[6] , \u_div/QInv[5] , 
        \u_div/QInv[4] , \u_div/QInv[3] , \u_div/QInv[2] , \u_div/QInv[1] , 
        \u_div/QInv[0] }), .sum(quotient) );
  MX2XL \u_div/u_mx_PartRem_1_2_0  ( .A(\u_div/PartRem[3][0] ), .B(
        \u_div/PartRem[3][0] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/SumTmp[1][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_0  ( .A(\u_div/PartRem[7][0] ), .B(
        \u_div/PartRem[7][0] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/SumTmp[5][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_5_1  ( .A(\u_div/SumTmp[5][1] ), .B(
        \u_div/SumTmp[5][1] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_0  ( .A(\u_div/PartRem[12][0] ), .B(
        \u_div/PartRem[12][0] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/SumTmp[10][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_0  ( .A(\u_div/PartRem[17][0] ), .B(
        \u_div/PartRem[17][0] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/SumTmp[15][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_15_1  ( .A(\u_div/SumTmp[15][1] ), .B(
        \u_div/SumTmp[15][1] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_0  ( .A(\u_div/PartRem[22][0] ), .B(
        \u_div/PartRem[22][0] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/SumTmp[20][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_20_1  ( .A(\u_div/SumTmp[20][1] ), .B(
        \u_div/SumTmp[20][1] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_0  ( .A(\u_div/PartRem[27][0] ), .B(
        \u_div/PartRem[27][0] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/SumTmp[25][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_25_1  ( .A(\u_div/SumTmp[25][1] ), .B(
        \u_div/SumTmp[25][1] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_0  ( .A(\u_div/PartRem[32][0] ), .B(
        \u_div/PartRem[32][0] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/SumTmp[30][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_30_1  ( .A(\u_div/SumTmp[30][1] ), .B(
        \u_div/SumTmp[30][1] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_0  ( .A(\u_div/PartRem[37][0] ), .B(
        \u_div/PartRem[37][0] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/SumTmp[35][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_35_1  ( .A(\u_div/SumTmp[35][1] ), .B(
        \u_div/SumTmp[35][1] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_0  ( .A(\u_div/PartRem[42][0] ), .B(
        \u_div/PartRem[42][0] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/SumTmp[40][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_40_1  ( .A(\u_div/SumTmp[40][1] ), .B(
        \u_div/SumTmp[40][1] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_0  ( .A(\u_div/PartRem[47][0] ), .B(
        \u_div/PartRem[47][0] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/SumTmp[45][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_45_1  ( .A(\u_div/SumTmp[45][1] ), .B(
        \u_div/SumTmp[45][1] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_0  ( .A(\u_div/PartRem[52][0] ), .B(
        \u_div/PartRem[52][0] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/SumTmp[50][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_50_1  ( .A(\u_div/SumTmp[50][1] ), .B(
        \u_div/SumTmp[50][1] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_55_1  ( .A(\u_div/SumTmp[55][1] ), .B(
        \u_div/SumTmp[55][1] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_0  ( .A(\u_div/PartRem[4][0] ), .B(
        \u_div/PartRem[4][0] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/SumTmp[2][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_0  ( .A(\u_div/PartRem[5][0] ), .B(
        \u_div/PartRem[5][0] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/SumTmp[3][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_0  ( .A(\u_div/PartRem[13][0] ), .B(
        \u_div/PartRem[13][0] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/SumTmp[11][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_0  ( .A(\u_div/PartRem[14][0] ), .B(
        \u_div/PartRem[14][0] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/SumTmp[12][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_0  ( .A(\u_div/PartRem[15][0] ), .B(
        \u_div/PartRem[15][0] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/SumTmp[13][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_0  ( .A(\u_div/PartRem[18][0] ), .B(
        \u_div/PartRem[18][0] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/SumTmp[16][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_0  ( .A(\u_div/PartRem[19][0] ), .B(
        \u_div/PartRem[19][0] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/SumTmp[17][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_0  ( .A(\u_div/PartRem[23][0] ), .B(
        \u_div/PartRem[23][0] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/SumTmp[21][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_0  ( .A(\u_div/PartRem[24][0] ), .B(
        \u_div/PartRem[24][0] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/SumTmp[22][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_0  ( .A(\u_div/PartRem[25][0] ), .B(
        \u_div/PartRem[25][0] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/SumTmp[23][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_0  ( .A(\u_div/PartRem[28][0] ), .B(
        \u_div/PartRem[28][0] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/SumTmp[26][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_0  ( .A(\u_div/PartRem[30][0] ), .B(
        \u_div/PartRem[30][0] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/SumTmp[28][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_0  ( .A(\u_div/PartRem[33][0] ), .B(
        \u_div/PartRem[33][0] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/SumTmp[31][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_0  ( .A(\u_div/PartRem[34][0] ), .B(
        \u_div/PartRem[34][0] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/SumTmp[32][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_0  ( .A(\u_div/PartRem[35][0] ), .B(
        \u_div/PartRem[35][0] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/SumTmp[33][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_0  ( .A(\u_div/PartRem[38][0] ), .B(
        \u_div/PartRem[38][0] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/SumTmp[36][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_0  ( .A(\u_div/PartRem[40][0] ), .B(
        \u_div/PartRem[40][0] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/SumTmp[38][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_0  ( .A(\u_div/PartRem[43][0] ), .B(
        \u_div/PartRem[43][0] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/SumTmp[41][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_0  ( .A(\u_div/PartRem[44][0] ), .B(
        \u_div/PartRem[44][0] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/SumTmp[42][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_0  ( .A(\u_div/PartRem[45][0] ), .B(
        \u_div/PartRem[45][0] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/SumTmp[43][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_0  ( .A(\u_div/PartRem[48][0] ), .B(
        \u_div/PartRem[48][0] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/SumTmp[46][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_0  ( .A(\u_div/PartRem[53][0] ), .B(
        \u_div/PartRem[53][0] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/SumTmp[51][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_0  ( .A(\u_div/PartRem[55][0] ), .B(
        \u_div/PartRem[55][0] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/SumTmp[53][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_0  ( .A(\u_div/PartRem[58][0] ), .B(
        \u_div/PartRem[58][0] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/SumTmp[56][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_0  ( .A(\u_div/PartRem[59][0] ), .B(
        \u_div/PartRem[59][0] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/SumTmp[57][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_0  ( .A(\u_div/PartRem[60][0] ), .B(
        \u_div/PartRem[60][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/SumTmp[58][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_59_1  ( .A(\u_div/PartRem[61][0] ), .B(
        \u_div/PartRem[61][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_1_3  ( .A(\u_div/PartRem[2][3] ), .B(
        \u_div/SumTmp[1][3] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_3  ( .A(\u_div/PartRem[3][3] ), .B(
        \u_div/SumTmp[2][3] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_3  ( .A(\u_div/PartRem[5][3] ), .B(
        \u_div/SumTmp[4][3] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_3  ( .A(\u_div/PartRem[7][3] ), .B(
        \u_div/SumTmp[6][3] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_9_3  ( .A(\u_div/PartRem[10][3] ), .B(
        \u_div/SumTmp[9][3] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_3  ( .A(\u_div/PartRem[12][3] ), .B(
        \u_div/SumTmp[11][3] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_3  ( .A(\u_div/PartRem[13][3] ), .B(
        \u_div/SumTmp[12][3] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_3  ( .A(\u_div/PartRem[15][3] ), .B(
        \u_div/SumTmp[14][3] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_3  ( .A(\u_div/PartRem[17][3] ), .B(
        \u_div/SumTmp[16][3] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_3  ( .A(\u_div/PartRem[18][3] ), .B(
        \u_div/SumTmp[17][3] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_3  ( .A(\u_div/PartRem[20][3] ), .B(
        \u_div/SumTmp[19][3] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_3  ( .A(\u_div/PartRem[22][3] ), .B(
        \u_div/SumTmp[21][3] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_3  ( .A(\u_div/PartRem[23][3] ), .B(
        \u_div/SumTmp[22][3] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_3  ( .A(\u_div/PartRem[25][3] ), .B(
        \u_div/SumTmp[24][3] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_3  ( .A(\u_div/PartRem[27][3] ), .B(
        \u_div/SumTmp[26][3] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_3  ( .A(\u_div/PartRem[28][3] ), .B(
        \u_div/SumTmp[27][3] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_3  ( .A(\u_div/PartRem[30][3] ), .B(
        \u_div/SumTmp[29][3] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_3  ( .A(\u_div/PartRem[32][3] ), .B(
        \u_div/SumTmp[31][3] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_3  ( .A(\u_div/PartRem[33][3] ), .B(
        \u_div/SumTmp[32][3] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_3  ( .A(\u_div/PartRem[35][3] ), .B(
        \u_div/SumTmp[34][3] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_3  ( .A(\u_div/PartRem[37][3] ), .B(
        \u_div/SumTmp[36][3] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_3  ( .A(\u_div/PartRem[38][3] ), .B(
        \u_div/SumTmp[37][3] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_3  ( .A(\u_div/PartRem[40][3] ), .B(
        \u_div/SumTmp[39][3] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_3  ( .A(\u_div/PartRem[42][3] ), .B(
        \u_div/SumTmp[41][3] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_3  ( .A(\u_div/PartRem[43][3] ), .B(
        \u_div/SumTmp[42][3] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_3  ( .A(\u_div/PartRem[45][3] ), .B(
        \u_div/SumTmp[44][3] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_3  ( .A(\u_div/PartRem[47][3] ), .B(
        \u_div/SumTmp[46][3] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_3  ( .A(\u_div/PartRem[48][3] ), .B(
        \u_div/SumTmp[47][3] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_3  ( .A(\u_div/PartRem[50][3] ), .B(
        \u_div/SumTmp[49][3] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_3  ( .A(\u_div/PartRem[52][3] ), .B(
        \u_div/SumTmp[51][3] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_3  ( .A(\u_div/PartRem[53][3] ), .B(
        \u_div/SumTmp[52][3] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_3  ( .A(\u_div/PartRem[55][3] ), .B(
        \u_div/SumTmp[54][3] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_3  ( .A(\u_div/PartRem[57][3] ), .B(
        \u_div/SumTmp[56][3] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_3  ( .A(\u_div/PartRem[58][3] ), .B(
        \u_div/SumTmp[57][3] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_3  ( .A(\u_div/PartRem[59][3] ), .B(
        \u_div/SumTmp[58][3] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_3  ( .A(\u_div/PartRem[63][0] ), .B(
        \u_div/SumTmp[59][3] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_3  ( .A(\u_div/PartRem[4][3] ), .B(
        \u_div/SumTmp[3][3] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_8_3  ( .A(\u_div/PartRem[9][3] ), .B(
        \u_div/SumTmp[8][3] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_3  ( .A(\u_div/PartRem[14][3] ), .B(
        \u_div/SumTmp[13][3] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_3  ( .A(\u_div/PartRem[19][3] ), .B(
        \u_div/SumTmp[18][3] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_3  ( .A(\u_div/PartRem[24][3] ), .B(
        \u_div/SumTmp[23][3] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_3  ( .A(\u_div/PartRem[29][3] ), .B(
        \u_div/SumTmp[28][3] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_3  ( .A(\u_div/PartRem[34][3] ), .B(
        \u_div/SumTmp[33][3] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_3  ( .A(\u_div/PartRem[39][3] ), .B(
        \u_div/SumTmp[38][3] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_3  ( .A(\u_div/PartRem[44][3] ), .B(
        \u_div/SumTmp[43][3] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_3  ( .A(\u_div/PartRem[49][3] ), .B(
        \u_div/SumTmp[48][3] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_3  ( .A(\u_div/PartRem[54][3] ), .B(
        \u_div/SumTmp[53][3] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/SumTmp[1][2] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][3] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_4  ( .A(\u_div/PartRem[64][0] ), .B(
        \u_div/SumTmp[59][4] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_3_1  ( .A(\u_div/SumTmp[3][1] ), .B(
        \u_div/SumTmp[3][1] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_4_1  ( .A(\u_div/SumTmp[4][1] ), .B(
        \u_div/SumTmp[4][1] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_0  ( .A(\u_div/PartRem[6][0] ), .B(
        \u_div/PartRem[6][0] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/SumTmp[4][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_13_1  ( .A(\u_div/SumTmp[13][1] ), .B(
        \u_div/SumTmp[13][1] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_18_1  ( .A(\u_div/SumTmp[18][1] ), .B(
        \u_div/SumTmp[18][1] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_0  ( .A(\u_div/PartRem[11][0] ), .B(
        \u_div/PartRem[11][0] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/SumTmp[9][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_14_1  ( .A(\u_div/SumTmp[14][1] ), .B(
        \u_div/SumTmp[14][1] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_0  ( .A(\u_div/PartRem[16][0] ), .B(
        \u_div/PartRem[16][0] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/SumTmp[14][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_0  ( .A(\u_div/PartRem[21][0] ), .B(
        \u_div/PartRem[21][0] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/SumTmp[19][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_12_1  ( .A(\u_div/SumTmp[12][1] ), .B(
        \u_div/SumTmp[12][1] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_17_1  ( .A(\u_div/SumTmp[17][1] ), .B(
        \u_div/SumTmp[17][1] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_6_1  ( .A(\u_div/SumTmp[6][1] ), .B(
        \u_div/SumTmp[6][1] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_22_1  ( .A(\u_div/SumTmp[22][1] ), .B(
        \u_div/SumTmp[22][1] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_11_1  ( .A(\u_div/SumTmp[11][1] ), .B(
        \u_div/SumTmp[11][1] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_16_1  ( .A(\u_div/SumTmp[16][1] ), .B(
        \u_div/SumTmp[16][1] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_23_1  ( .A(\u_div/SumTmp[23][1] ), .B(
        \u_div/SumTmp[23][1] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_21_1  ( .A(\u_div/SumTmp[21][1] ), .B(
        \u_div/SumTmp[21][1] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_24_1  ( .A(\u_div/SumTmp[24][1] ), .B(
        \u_div/SumTmp[24][1] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_0  ( .A(\u_div/PartRem[26][0] ), .B(
        \u_div/PartRem[26][0] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/SumTmp[24][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_26_1  ( .A(\u_div/SumTmp[26][1] ), .B(
        \u_div/SumTmp[26][1] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_27_1  ( .A(\u_div/SumTmp[27][1] ), .B(
        \u_div/SumTmp[27][1] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_29_1  ( .A(\u_div/SumTmp[29][1] ), .B(
        \u_div/SumTmp[29][1] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_0  ( .A(\u_div/PartRem[31][0] ), .B(
        \u_div/PartRem[31][0] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/SumTmp[29][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_31_1  ( .A(\u_div/SumTmp[31][1] ), .B(
        \u_div/SumTmp[31][1] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_32_1  ( .A(\u_div/SumTmp[32][1] ), .B(
        \u_div/SumTmp[32][1] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_33_1  ( .A(\u_div/SumTmp[33][1] ), .B(
        \u_div/SumTmp[33][1] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_34_1  ( .A(\u_div/SumTmp[34][1] ), .B(
        \u_div/SumTmp[34][1] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_0  ( .A(\u_div/PartRem[36][0] ), .B(
        \u_div/PartRem[36][0] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/SumTmp[34][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_36_1  ( .A(\u_div/SumTmp[36][1] ), .B(
        \u_div/SumTmp[36][1] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_37_1  ( .A(\u_div/SumTmp[37][1] ), .B(
        \u_div/SumTmp[37][1] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_39_1  ( .A(\u_div/SumTmp[39][1] ), .B(
        \u_div/SumTmp[39][1] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_0  ( .A(\u_div/PartRem[41][0] ), .B(
        \u_div/PartRem[41][0] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/SumTmp[39][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_41_1  ( .A(\u_div/SumTmp[41][1] ), .B(
        \u_div/SumTmp[41][1] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_42_1  ( .A(\u_div/SumTmp[42][1] ), .B(
        \u_div/SumTmp[42][1] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_43_1  ( .A(\u_div/SumTmp[43][1] ), .B(
        \u_div/SumTmp[43][1] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_44_1  ( .A(\u_div/SumTmp[44][1] ), .B(
        \u_div/SumTmp[44][1] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_0  ( .A(\u_div/PartRem[46][0] ), .B(
        \u_div/PartRem[46][0] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/SumTmp[44][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_46_1  ( .A(\u_div/SumTmp[46][1] ), .B(
        \u_div/SumTmp[46][1] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_47_1  ( .A(\u_div/SumTmp[47][1] ), .B(
        \u_div/SumTmp[47][1] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_0  ( .A(\u_div/PartRem[51][0] ), .B(
        \u_div/PartRem[51][0] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/SumTmp[49][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_51_1  ( .A(\u_div/SumTmp[51][1] ), .B(
        \u_div/SumTmp[51][1] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_52_1  ( .A(\u_div/SumTmp[52][1] ), .B(
        \u_div/SumTmp[52][1] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_54_1  ( .A(\u_div/SumTmp[54][1] ), .B(
        \u_div/SumTmp[54][1] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_0  ( .A(\u_div/PartRem[56][0] ), .B(
        \u_div/PartRem[56][0] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/SumTmp[54][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_57_1  ( .A(\u_div/SumTmp[57][1] ), .B(
        \u_div/SumTmp[57][1] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_58_1  ( .A(\u_div/SumTmp[58][1] ), .B(
        \u_div/SumTmp[58][1] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_2_1  ( .A(\u_div/SumTmp[2][1] ), .B(
        \u_div/SumTmp[2][1] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_3  ( .A(\u_div/PartRem[6][3] ), .B(
        \u_div/SumTmp[5][3] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_3  ( .A(\u_div/PartRem[11][3] ), .B(
        \u_div/SumTmp[10][3] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_3  ( .A(\u_div/PartRem[16][3] ), .B(
        \u_div/SumTmp[15][3] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_3  ( .A(\u_div/PartRem[21][3] ), .B(
        \u_div/SumTmp[20][3] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_3  ( .A(\u_div/PartRem[26][3] ), .B(
        \u_div/SumTmp[25][3] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_3  ( .A(\u_div/PartRem[31][3] ), .B(
        \u_div/SumTmp[30][3] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_3  ( .A(\u_div/PartRem[36][3] ), .B(
        \u_div/SumTmp[35][3] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_3  ( .A(\u_div/PartRem[41][3] ), .B(
        \u_div/SumTmp[40][3] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_3  ( .A(\u_div/PartRem[46][3] ), .B(
        \u_div/SumTmp[45][3] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_3  ( .A(\u_div/PartRem[51][3] ), .B(
        \u_div/SumTmp[50][3] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_3  ( .A(\u_div/PartRem[56][3] ), .B(
        \u_div/SumTmp[55][3] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_1_4  ( .A(\u_div/PartRem[2][4] ), .B(
        \u_div/SumTmp[1][4] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_4  ( .A(\u_div/PartRem[7][4] ), .B(
        \u_div/SumTmp[6][4] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_4  ( .A(\u_div/PartRem[12][4] ), .B(
        \u_div/SumTmp[11][4] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_4  ( .A(\u_div/PartRem[17][4] ), .B(
        \u_div/SumTmp[16][4] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_4  ( .A(\u_div/PartRem[22][4] ), .B(
        \u_div/SumTmp[21][4] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_4  ( .A(\u_div/PartRem[27][4] ), .B(
        \u_div/SumTmp[26][4] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_4  ( .A(\u_div/PartRem[32][4] ), .B(
        \u_div/SumTmp[31][4] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_4  ( .A(\u_div/PartRem[37][4] ), .B(
        \u_div/SumTmp[36][4] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_4  ( .A(\u_div/PartRem[42][4] ), .B(
        \u_div/SumTmp[41][4] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_4  ( .A(\u_div/PartRem[47][4] ), .B(
        \u_div/SumTmp[46][4] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_4  ( .A(\u_div/PartRem[52][4] ), .B(
        \u_div/SumTmp[51][4] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_4  ( .A(\u_div/PartRem[3][4] ), .B(
        \u_div/SumTmp[2][4] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_4  ( .A(\u_div/PartRem[4][4] ), .B(
        \u_div/SumTmp[3][4] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_4  ( .A(\u_div/PartRem[5][4] ), .B(
        \u_div/SumTmp[4][4] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_4  ( .A(\u_div/PartRem[6][4] ), .B(
        \u_div/SumTmp[5][4] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_4  ( .A(\u_div/PartRem[8][4] ), .B(
        \u_div/SumTmp[7][4] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_4  ( .A(\u_div/PartRem[15][4] ), .B(
        \u_div/SumTmp[14][4] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_4  ( .A(\u_div/PartRem[14][4] ), .B(
        \u_div/SumTmp[13][4] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_4  ( .A(\u_div/PartRem[19][4] ), .B(
        \u_div/SumTmp[18][4] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_4  ( .A(\u_div/PartRem[13][4] ), .B(
        \u_div/SumTmp[12][4] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_4  ( .A(\u_div/PartRem[18][4] ), .B(
        \u_div/SumTmp[17][4] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_4  ( .A(\u_div/PartRem[11][4] ), .B(
        \u_div/SumTmp[10][4] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_4  ( .A(\u_div/PartRem[16][4] ), .B(
        \u_div/SumTmp[15][4] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_4  ( .A(\u_div/PartRem[21][4] ), .B(
        \u_div/SumTmp[20][4] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_4  ( .A(\u_div/PartRem[23][4] ), .B(
        \u_div/SumTmp[22][4] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_4  ( .A(\u_div/PartRem[26][4] ), .B(
        \u_div/SumTmp[25][4] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_4  ( .A(\u_div/PartRem[24][4] ), .B(
        \u_div/SumTmp[23][4] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_4  ( .A(\u_div/PartRem[25][4] ), .B(
        \u_div/SumTmp[24][4] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_4  ( .A(\u_div/PartRem[28][4] ), .B(
        \u_div/SumTmp[27][4] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_4  ( .A(\u_div/PartRem[30][4] ), .B(
        \u_div/SumTmp[29][4] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_4  ( .A(\u_div/PartRem[31][4] ), .B(
        \u_div/SumTmp[30][4] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_4  ( .A(\u_div/PartRem[34][4] ), .B(
        \u_div/SumTmp[33][4] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_4  ( .A(\u_div/PartRem[33][4] ), .B(
        \u_div/SumTmp[32][4] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_4  ( .A(\u_div/PartRem[35][4] ), .B(
        \u_div/SumTmp[34][4] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_4  ( .A(\u_div/PartRem[36][4] ), .B(
        \u_div/SumTmp[35][4] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_4  ( .A(\u_div/PartRem[38][4] ), .B(
        \u_div/SumTmp[37][4] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_4  ( .A(\u_div/PartRem[40][4] ), .B(
        \u_div/SumTmp[39][4] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_4  ( .A(\u_div/PartRem[41][4] ), .B(
        \u_div/SumTmp[40][4] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_4  ( .A(\u_div/PartRem[44][4] ), .B(
        \u_div/SumTmp[43][4] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_4  ( .A(\u_div/PartRem[43][4] ), .B(
        \u_div/SumTmp[42][4] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_4  ( .A(\u_div/PartRem[45][4] ), .B(
        \u_div/SumTmp[44][4] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_4  ( .A(\u_div/PartRem[46][4] ), .B(
        \u_div/SumTmp[45][4] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_4  ( .A(\u_div/PartRem[48][4] ), .B(
        \u_div/SumTmp[47][4] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_4  ( .A(\u_div/PartRem[51][4] ), .B(
        \u_div/SumTmp[50][4] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_4  ( .A(\u_div/PartRem[55][4] ), .B(
        \u_div/SumTmp[54][4] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_4  ( .A(\u_div/PartRem[53][4] ), .B(
        \u_div/SumTmp[52][4] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_4  ( .A(\u_div/PartRem[58][4] ), .B(
        \u_div/SumTmp[57][4] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_4  ( .A(\u_div/PartRem[56][4] ), .B(
        \u_div/SumTmp[55][4] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_4  ( .A(\u_div/PartRem[59][4] ), .B(
        \u_div/SumTmp[58][4] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_8_4  ( .A(\u_div/PartRem[9][4] ), .B(
        \u_div/SumTmp[8][4] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][5] ) );
  CLKMX2X6 \u_div/u_mx_PartRem_1_8_1  ( .A(\u_div/SumTmp[8][1] ), .B(
        \u_div/SumTmp[8][1] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_8_0  ( .A(\u_div/PartRem[9][0] ), .B(
        \u_div/PartRem[9][0] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/SumTmp[7][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_9_4  ( .A(\u_div/PartRem[10][4] ), .B(
        \u_div/SumTmp[9][4] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][5] ) );
  MX2X6 \u_div/u_mx_PartRem_1_9_1  ( .A(\u_div/SumTmp[9][1] ), .B(
        \u_div/SumTmp[9][1] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_9_0  ( .A(\u_div/PartRem[10][0] ), .B(
        \u_div/PartRem[10][0] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/SumTmp[8][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_19_4  ( .A(\u_div/PartRem[20][4] ), .B(
        \u_div/SumTmp[19][4] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][5] ) );
  MX2X6 \u_div/u_mx_PartRem_1_19_1  ( .A(\u_div/SumTmp[19][1] ), .B(
        \u_div/SumTmp[19][1] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_19_0  ( .A(\u_div/PartRem[20][0] ), .B(
        \u_div/PartRem[20][0] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/SumTmp[18][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_28_4  ( .A(\u_div/PartRem[29][4] ), .B(
        \u_div/SumTmp[28][4] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][5] ) );
  CLKMX2X6 \u_div/u_mx_PartRem_1_28_1  ( .A(\u_div/SumTmp[28][1] ), .B(
        \u_div/SumTmp[28][1] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_28_0  ( .A(\u_div/PartRem[29][0] ), .B(
        \u_div/PartRem[29][0] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/SumTmp[27][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_38_4  ( .A(\u_div/PartRem[39][4] ), .B(
        \u_div/SumTmp[38][4] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][5] ) );
  CLKMX2X6 \u_div/u_mx_PartRem_1_38_1  ( .A(\u_div/SumTmp[38][1] ), .B(
        \u_div/SumTmp[38][1] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_38_0  ( .A(\u_div/PartRem[39][0] ), .B(
        \u_div/PartRem[39][0] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/SumTmp[37][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_48_4  ( .A(\u_div/PartRem[49][4] ), .B(
        \u_div/SumTmp[48][4] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][5] ) );
  CLKMX2X6 \u_div/u_mx_PartRem_1_48_1  ( .A(\u_div/SumTmp[48][1] ), .B(
        \u_div/SumTmp[48][1] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_48_0  ( .A(\u_div/PartRem[49][0] ), .B(
        \u_div/PartRem[49][0] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/SumTmp[47][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_49_4  ( .A(\u_div/PartRem[50][4] ), .B(
        \u_div/SumTmp[49][4] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][5] ) );
  MX2X6 \u_div/u_mx_PartRem_1_49_1  ( .A(\u_div/SumTmp[49][1] ), .B(
        \u_div/SumTmp[49][1] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_49_0  ( .A(\u_div/PartRem[50][0] ), .B(
        \u_div/PartRem[50][0] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/SumTmp[48][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_53_4  ( .A(\u_div/PartRem[54][4] ), .B(
        \u_div/SumTmp[53][4] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][5] ) );
  CLKMX2X6 \u_div/u_mx_PartRem_1_53_1  ( .A(\u_div/SumTmp[53][1] ), .B(
        \u_div/SumTmp[53][1] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_53_0  ( .A(\u_div/PartRem[54][0] ), .B(
        \u_div/PartRem[54][0] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/SumTmp[52][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_56_4  ( .A(\u_div/PartRem[57][4] ), .B(
        \u_div/SumTmp[56][4] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][5] ) );
  CLKMX2X6 \u_div/u_mx_PartRem_1_56_1  ( .A(\u_div/SumTmp[56][1] ), .B(
        \u_div/SumTmp[56][1] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_56_0  ( .A(\u_div/PartRem[57][0] ), .B(
        \u_div/PartRem[57][0] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/SumTmp[55][1] ) );
  MX2X6 \u_div/u_mx_PartRem_1_7_1  ( .A(\u_div/SumTmp[7][1] ), .B(
        \u_div/SumTmp[7][1] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][2] ) );
  MX2X4 \u_div/u_mx_PartRem_1_7_3  ( .A(\u_div/PartRem[8][3] ), .B(
        \u_div/SumTmp[7][3] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][4] ) );
  MX2X1 \u_div/u_mx_PartRem_1_7_0  ( .A(\u_div/PartRem[8][0] ), .B(
        \u_div/PartRem[8][0] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/SumTmp[6][1] ) );
  CLKMX2X8 \u_div/u_mx_PartRem_1_10_1  ( .A(\u_div/SumTmp[10][1] ), .B(
        \u_div/SumTmp[10][1] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][2] ) );
  OR2X6 U1 ( .A(\u_div/PartRem[11][5] ), .B(\u_div/u_add_PartRem_2_10/n2 ), 
        .Y(\u_div/CryTmp[10][6] ) );
  MXI2X4 U2 ( .A(\u_div/SumTmp[7][2] ), .B(\u_div/PartRem[8][2] ), .S0(
        \u_div/CryTmp[7][6] ), .Y(\u_div/PartRem[7][3] ) );
  OR2X6 U3 ( .A(\u_div/PartRem[8][5] ), .B(\u_div/u_add_PartRem_2_7/n2 ), .Y(
        \u_div/CryTmp[7][6] ) );
  OR2X8 U4 ( .A(\u_div/PartRem[7][5] ), .B(\u_div/u_add_PartRem_2_6/n2 ), .Y(
        \u_div/CryTmp[6][6] ) );
  ADDHX2 U5 ( .A(\u_div/PartRem[7][4] ), .B(\u_div/u_add_PartRem_2_6/n3 ), 
        .CO(\u_div/u_add_PartRem_2_6/n2 ), .S(\u_div/SumTmp[6][4] ) );
  OR2X8 U6 ( .A(\u_div/PartRem[6][5] ), .B(\u_div/u_add_PartRem_2_5/n2 ), .Y(
        \u_div/CryTmp[5][6] ) );
  ADDHX2 U7 ( .A(\u_div/PartRem[6][4] ), .B(\u_div/u_add_PartRem_2_5/n3 ), 
        .CO(\u_div/u_add_PartRem_2_5/n2 ), .S(\u_div/SumTmp[5][4] ) );
  OR2X8 U8 ( .A(\u_div/PartRem[5][5] ), .B(\u_div/u_add_PartRem_2_4/n2 ), .Y(
        \u_div/CryTmp[4][6] ) );
  ADDHX2 U9 ( .A(\u_div/PartRem[5][4] ), .B(\u_div/u_add_PartRem_2_4/n3 ), 
        .CO(\u_div/u_add_PartRem_2_4/n2 ), .S(\u_div/SumTmp[4][4] ) );
  OR2X8 U10 ( .A(\u_div/PartRem[4][5] ), .B(\u_div/u_add_PartRem_2_3/n2 ), .Y(
        \u_div/CryTmp[3][6] ) );
  ADDHX2 U11 ( .A(\u_div/PartRem[4][4] ), .B(\u_div/u_add_PartRem_2_3/n3 ), 
        .CO(\u_div/u_add_PartRem_2_3/n2 ), .S(\u_div/SumTmp[3][4] ) );
  OR2X8 U12 ( .A(\u_div/PartRem[3][5] ), .B(\u_div/u_add_PartRem_2_2/n2 ), .Y(
        \u_div/CryTmp[2][6] ) );
  ADDHX2 U13 ( .A(\u_div/PartRem[3][4] ), .B(\u_div/u_add_PartRem_2_2/n3 ), 
        .CO(\u_div/u_add_PartRem_2_2/n2 ), .S(\u_div/SumTmp[2][4] ) );
  OR2X8 U14 ( .A(\u_div/PartRem[59][5] ), .B(\u_div/u_add_PartRem_2_58/n2 ), 
        .Y(\u_div/CryTmp[58][6] ) );
  ADDHX2 U15 ( .A(\u_div/PartRem[59][4] ), .B(\u_div/u_add_PartRem_2_58/n3 ), 
        .CO(\u_div/u_add_PartRem_2_58/n2 ), .S(\u_div/SumTmp[58][4] ) );
  XOR2XL U16 ( .A(\u_div/CryTmp[56][6] ), .B(n3), .Y(\u_div/QInv[56] ) );
  MXI2X4 U17 ( .A(\u_div/SumTmp[56][2] ), .B(\u_div/PartRem[57][2] ), .S0(
        \u_div/CryTmp[56][6] ), .Y(\u_div/PartRem[56][3] ) );
  OR2X6 U18 ( .A(\u_div/PartRem[57][5] ), .B(\u_div/u_add_PartRem_2_56/n2 ), 
        .Y(\u_div/CryTmp[56][6] ) );
  XOR2XL U19 ( .A(\u_div/CryTmp[53][6] ), .B(n3), .Y(\u_div/QInv[53] ) );
  MXI2X4 U20 ( .A(\u_div/SumTmp[53][2] ), .B(\u_div/PartRem[54][2] ), .S0(
        \u_div/CryTmp[53][6] ), .Y(\u_div/PartRem[53][3] ) );
  OR2X6 U21 ( .A(\u_div/PartRem[54][5] ), .B(\u_div/u_add_PartRem_2_53/n2 ), 
        .Y(\u_div/CryTmp[53][6] ) );
  XOR2XL U22 ( .A(\u_div/CryTmp[49][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[49] ) );
  MXI2X4 U23 ( .A(\u_div/SumTmp[49][2] ), .B(\u_div/PartRem[50][2] ), .S0(
        \u_div/CryTmp[49][6] ), .Y(\u_div/PartRem[49][3] ) );
  OR2X6 U24 ( .A(\u_div/PartRem[50][5] ), .B(\u_div/u_add_PartRem_2_49/n2 ), 
        .Y(\u_div/CryTmp[49][6] ) );
  XOR2XL U25 ( .A(\u_div/CryTmp[48][6] ), .B(n3), .Y(\u_div/QInv[48] ) );
  MXI2X4 U26 ( .A(\u_div/SumTmp[48][2] ), .B(\u_div/PartRem[49][2] ), .S0(
        \u_div/CryTmp[48][6] ), .Y(\u_div/PartRem[48][3] ) );
  OR2X6 U27 ( .A(\u_div/PartRem[49][5] ), .B(\u_div/u_add_PartRem_2_48/n2 ), 
        .Y(\u_div/CryTmp[48][6] ) );
  OR2X8 U28 ( .A(\u_div/PartRem[40][5] ), .B(\u_div/u_add_PartRem_2_39/n2 ), 
        .Y(\u_div/CryTmp[39][6] ) );
  ADDHX2 U29 ( .A(\u_div/PartRem[40][4] ), .B(\u_div/u_add_PartRem_2_39/n3 ), 
        .CO(\u_div/u_add_PartRem_2_39/n2 ), .S(\u_div/SumTmp[39][4] ) );
  XOR2XL U30 ( .A(\u_div/CryTmp[38][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[38] ) );
  MXI2X4 U31 ( .A(\u_div/SumTmp[38][2] ), .B(\u_div/PartRem[39][2] ), .S0(
        \u_div/CryTmp[38][6] ), .Y(\u_div/PartRem[38][3] ) );
  OR2X6 U32 ( .A(\u_div/PartRem[39][5] ), .B(\u_div/u_add_PartRem_2_38/n2 ), 
        .Y(\u_div/CryTmp[38][6] ) );
  OR2X8 U33 ( .A(\u_div/PartRem[30][5] ), .B(\u_div/u_add_PartRem_2_29/n2 ), 
        .Y(\u_div/CryTmp[29][6] ) );
  ADDHX2 U34 ( .A(\u_div/PartRem[30][4] ), .B(\u_div/u_add_PartRem_2_29/n3 ), 
        .CO(\u_div/u_add_PartRem_2_29/n2 ), .S(\u_div/SumTmp[29][4] ) );
  XOR2XL U35 ( .A(\u_div/CryTmp[28][6] ), .B(n5), .Y(\u_div/QInv[28] ) );
  MXI2X4 U36 ( .A(\u_div/SumTmp[28][2] ), .B(\u_div/PartRem[29][2] ), .S0(
        \u_div/CryTmp[28][6] ), .Y(\u_div/PartRem[28][3] ) );
  OR2X6 U37 ( .A(\u_div/PartRem[29][5] ), .B(\u_div/u_add_PartRem_2_28/n2 ), 
        .Y(\u_div/CryTmp[28][6] ) );
  XOR2XL U38 ( .A(\u_div/CryTmp[19][6] ), .B(n3), .Y(\u_div/QInv[19] ) );
  MXI2X4 U39 ( .A(\u_div/SumTmp[19][2] ), .B(\u_div/PartRem[20][2] ), .S0(
        \u_div/CryTmp[19][6] ), .Y(\u_div/PartRem[19][3] ) );
  OR2X6 U40 ( .A(\u_div/PartRem[20][5] ), .B(\u_div/u_add_PartRem_2_19/n2 ), 
        .Y(\u_div/CryTmp[19][6] ) );
  OR2X8 U41 ( .A(\u_div/PartRem[19][5] ), .B(\u_div/u_add_PartRem_2_18/n2 ), 
        .Y(\u_div/CryTmp[18][6] ) );
  ADDHX2 U42 ( .A(\u_div/PartRem[19][4] ), .B(\u_div/u_add_PartRem_2_18/n3 ), 
        .CO(\u_div/u_add_PartRem_2_18/n2 ), .S(\u_div/SumTmp[18][4] ) );
  XOR2XL U43 ( .A(\u_div/CryTmp[9][6] ), .B(n3), .Y(\u_div/QInv[9] ) );
  MXI2X4 U44 ( .A(\u_div/SumTmp[9][2] ), .B(\u_div/PartRem[10][2] ), .S0(
        \u_div/CryTmp[9][6] ), .Y(\u_div/PartRem[9][3] ) );
  OR2X6 U45 ( .A(\u_div/PartRem[10][5] ), .B(\u_div/u_add_PartRem_2_9/n2 ), 
        .Y(\u_div/CryTmp[9][6] ) );
  XOR2XL U46 ( .A(\u_div/CryTmp[8][6] ), .B(n3), .Y(\u_div/QInv[8] ) );
  MXI2X4 U47 ( .A(\u_div/SumTmp[8][2] ), .B(\u_div/PartRem[9][2] ), .S0(
        \u_div/CryTmp[8][6] ), .Y(\u_div/PartRem[8][3] ) );
  OR2X6 U48 ( .A(\u_div/PartRem[9][5] ), .B(\u_div/u_add_PartRem_2_8/n2 ), .Y(
        \u_div/CryTmp[8][6] ) );
  MXI2X1 U49 ( .A(\u_div/SumTmp[13][2] ), .B(\u_div/PartRem[14][2] ), .S0(
        \u_div/CryTmp[13][6] ), .Y(\u_div/PartRem[13][3] ) );
  MXI2X1 U50 ( .A(\u_div/SumTmp[18][2] ), .B(\u_div/PartRem[19][2] ), .S0(
        \u_div/CryTmp[18][6] ), .Y(\u_div/PartRem[18][3] ) );
  MXI2X1 U51 ( .A(\u_div/SumTmp[23][2] ), .B(\u_div/PartRem[24][2] ), .S0(
        \u_div/CryTmp[23][6] ), .Y(\u_div/PartRem[23][3] ) );
  MXI2X1 U52 ( .A(\u_div/SumTmp[33][2] ), .B(\u_div/PartRem[34][2] ), .S0(
        \u_div/CryTmp[33][6] ), .Y(\u_div/PartRem[33][3] ) );
  MXI2X1 U53 ( .A(\u_div/SumTmp[43][2] ), .B(\u_div/PartRem[44][2] ), .S0(
        \u_div/CryTmp[43][6] ), .Y(\u_div/PartRem[43][3] ) );
  ADDHXL U54 ( .A(\u_div/PartRem[13][4] ), .B(\u_div/u_add_PartRem_2_12/n3 ), 
        .CO(\u_div/u_add_PartRem_2_12/n2 ), .S(\u_div/SumTmp[12][4] ) );
  ADDHXL U55 ( .A(\u_div/PartRem[12][4] ), .B(\u_div/u_add_PartRem_2_11/n3 ), 
        .CO(\u_div/u_add_PartRem_2_11/n2 ), .S(\u_div/SumTmp[11][4] ) );
  OR2X1 U56 ( .A(\u_div/PartRem[12][2] ), .B(\u_div/PartRem[12][3] ), .Y(
        \u_div/u_add_PartRem_2_11/n3 ) );
  ADDHXL U57 ( .A(\u_div/PartRem[15][4] ), .B(\u_div/u_add_PartRem_2_14/n3 ), 
        .CO(\u_div/u_add_PartRem_2_14/n2 ), .S(\u_div/SumTmp[14][4] ) );
  OR2X1 U58 ( .A(\u_div/PartRem[15][2] ), .B(\u_div/PartRem[15][3] ), .Y(
        \u_div/u_add_PartRem_2_14/n3 ) );
  ADDHXL U59 ( .A(\u_div/PartRem[14][4] ), .B(\u_div/u_add_PartRem_2_13/n3 ), 
        .CO(\u_div/u_add_PartRem_2_13/n2 ), .S(\u_div/SumTmp[13][4] ) );
  OR2X1 U60 ( .A(\u_div/PartRem[14][2] ), .B(\u_div/PartRem[14][3] ), .Y(
        \u_div/u_add_PartRem_2_13/n3 ) );
  ADDHXL U61 ( .A(\u_div/PartRem[16][4] ), .B(\u_div/u_add_PartRem_2_15/n3 ), 
        .CO(\u_div/u_add_PartRem_2_15/n2 ), .S(\u_div/SumTmp[15][4] ) );
  OR2X1 U62 ( .A(\u_div/PartRem[16][2] ), .B(\u_div/PartRem[16][3] ), .Y(
        \u_div/u_add_PartRem_2_15/n3 ) );
  ADDHXL U63 ( .A(\u_div/PartRem[17][4] ), .B(\u_div/u_add_PartRem_2_16/n3 ), 
        .CO(\u_div/u_add_PartRem_2_16/n2 ), .S(\u_div/SumTmp[16][4] ) );
  OR2X1 U64 ( .A(\u_div/PartRem[17][2] ), .B(\u_div/PartRem[17][3] ), .Y(
        \u_div/u_add_PartRem_2_16/n3 ) );
  ADDHXL U65 ( .A(\u_div/PartRem[18][4] ), .B(\u_div/u_add_PartRem_2_17/n3 ), 
        .CO(\u_div/u_add_PartRem_2_17/n2 ), .S(\u_div/SumTmp[17][4] ) );
  OR2X1 U66 ( .A(\u_div/PartRem[19][2] ), .B(\u_div/PartRem[19][3] ), .Y(
        \u_div/u_add_PartRem_2_18/n3 ) );
  ADDHXL U67 ( .A(\u_div/PartRem[20][4] ), .B(\u_div/u_add_PartRem_2_19/n3 ), 
        .CO(\u_div/u_add_PartRem_2_19/n2 ), .S(\u_div/SumTmp[19][4] ) );
  OR2X1 U68 ( .A(\u_div/PartRem[20][2] ), .B(\u_div/PartRem[20][3] ), .Y(
        \u_div/u_add_PartRem_2_19/n3 ) );
  ADDHXL U69 ( .A(\u_div/PartRem[24][4] ), .B(\u_div/u_add_PartRem_2_23/n3 ), 
        .CO(\u_div/u_add_PartRem_2_23/n2 ), .S(\u_div/SumTmp[23][4] ) );
  OR2X1 U70 ( .A(\u_div/PartRem[24][2] ), .B(\u_div/PartRem[24][3] ), .Y(
        \u_div/u_add_PartRem_2_23/n3 ) );
  ADDHXL U71 ( .A(\u_div/PartRem[23][4] ), .B(\u_div/u_add_PartRem_2_22/n3 ), 
        .CO(\u_div/u_add_PartRem_2_22/n2 ), .S(\u_div/SumTmp[22][4] ) );
  ADDHXL U72 ( .A(\u_div/PartRem[22][4] ), .B(\u_div/u_add_PartRem_2_21/n3 ), 
        .CO(\u_div/u_add_PartRem_2_21/n2 ), .S(\u_div/SumTmp[21][4] ) );
  OR2X1 U73 ( .A(\u_div/PartRem[22][2] ), .B(\u_div/PartRem[22][3] ), .Y(
        \u_div/u_add_PartRem_2_21/n3 ) );
  ADDHXL U74 ( .A(\u_div/PartRem[21][4] ), .B(\u_div/u_add_PartRem_2_20/n3 ), 
        .CO(\u_div/u_add_PartRem_2_20/n2 ), .S(\u_div/SumTmp[20][4] ) );
  OR2X1 U75 ( .A(\u_div/PartRem[21][2] ), .B(\u_div/PartRem[21][3] ), .Y(
        \u_div/u_add_PartRem_2_20/n3 ) );
  MXI2X1 U76 ( .A(\u_div/SumTmp[3][2] ), .B(\u_div/PartRem[4][2] ), .S0(
        \u_div/CryTmp[3][6] ), .Y(\u_div/PartRem[3][3] ) );
  OR2X1 U77 ( .A(\u_div/PartRem[7][2] ), .B(\u_div/PartRem[7][3] ), .Y(
        \u_div/u_add_PartRem_2_6/n3 ) );
  ADDHXL U78 ( .A(\u_div/PartRem[11][4] ), .B(\u_div/u_add_PartRem_2_10/n3 ), 
        .CO(\u_div/u_add_PartRem_2_10/n2 ), .S(\u_div/SumTmp[10][4] ) );
  OR2X1 U79 ( .A(\u_div/PartRem[11][2] ), .B(\u_div/PartRem[11][3] ), .Y(
        \u_div/u_add_PartRem_2_10/n3 ) );
  OR2X1 U80 ( .A(\u_div/PartRem[4][2] ), .B(\u_div/PartRem[4][3] ), .Y(
        \u_div/u_add_PartRem_2_3/n3 ) );
  ADDHXL U81 ( .A(\u_div/PartRem[8][4] ), .B(\u_div/u_add_PartRem_2_7/n3 ), 
        .CO(\u_div/u_add_PartRem_2_7/n2 ), .S(\u_div/SumTmp[7][4] ) );
  ADDHXL U82 ( .A(\u_div/PartRem[10][4] ), .B(\u_div/u_add_PartRem_2_9/n3 ), 
        .CO(\u_div/u_add_PartRem_2_9/n2 ), .S(\u_div/SumTmp[9][4] ) );
  OR2X1 U83 ( .A(\u_div/PartRem[10][2] ), .B(\u_div/PartRem[10][3] ), .Y(
        \u_div/u_add_PartRem_2_9/n3 ) );
  ADDHXL U84 ( .A(\u_div/PartRem[9][4] ), .B(\u_div/u_add_PartRem_2_8/n3 ), 
        .CO(\u_div/u_add_PartRem_2_8/n2 ), .S(\u_div/SumTmp[8][4] ) );
  OR2X1 U85 ( .A(\u_div/PartRem[9][2] ), .B(\u_div/PartRem[9][3] ), .Y(
        \u_div/u_add_PartRem_2_8/n3 ) );
  OR2X1 U86 ( .A(\u_div/PartRem[6][2] ), .B(\u_div/PartRem[6][3] ), .Y(
        \u_div/u_add_PartRem_2_5/n3 ) );
  OR2X1 U87 ( .A(\u_div/PartRem[5][2] ), .B(\u_div/PartRem[5][3] ), .Y(
        \u_div/u_add_PartRem_2_4/n3 ) );
  ADDHXL U88 ( .A(\u_div/PartRem[25][4] ), .B(\u_div/u_add_PartRem_2_24/n3 ), 
        .CO(\u_div/u_add_PartRem_2_24/n2 ), .S(\u_div/SumTmp[24][4] ) );
  OR2X1 U89 ( .A(\u_div/PartRem[25][2] ), .B(\u_div/PartRem[25][3] ), .Y(
        \u_div/u_add_PartRem_2_24/n3 ) );
  ADDHXL U90 ( .A(\u_div/PartRem[26][4] ), .B(\u_div/u_add_PartRem_2_25/n3 ), 
        .CO(\u_div/u_add_PartRem_2_25/n2 ), .S(\u_div/SumTmp[25][4] ) );
  OR2X1 U91 ( .A(\u_div/PartRem[26][2] ), .B(\u_div/PartRem[26][3] ), .Y(
        \u_div/u_add_PartRem_2_25/n3 ) );
  ADDHXL U92 ( .A(\u_div/PartRem[27][4] ), .B(\u_div/u_add_PartRem_2_26/n3 ), 
        .CO(\u_div/u_add_PartRem_2_26/n2 ), .S(\u_div/SumTmp[26][4] ) );
  OR2X1 U93 ( .A(\u_div/PartRem[27][2] ), .B(\u_div/PartRem[27][3] ), .Y(
        \u_div/u_add_PartRem_2_26/n3 ) );
  ADDHXL U94 ( .A(\u_div/PartRem[28][4] ), .B(\u_div/u_add_PartRem_2_27/n3 ), 
        .CO(\u_div/u_add_PartRem_2_27/n2 ), .S(\u_div/SumTmp[27][4] ) );
  ADDHXL U95 ( .A(\u_div/PartRem[29][4] ), .B(\u_div/u_add_PartRem_2_28/n3 ), 
        .CO(\u_div/u_add_PartRem_2_28/n2 ), .S(\u_div/SumTmp[28][4] ) );
  OR2X1 U96 ( .A(\u_div/PartRem[29][2] ), .B(\u_div/PartRem[29][3] ), .Y(
        \u_div/u_add_PartRem_2_28/n3 ) );
  OR2X1 U97 ( .A(\u_div/PartRem[30][2] ), .B(\u_div/PartRem[30][3] ), .Y(
        \u_div/u_add_PartRem_2_29/n3 ) );
  ADDHXL U98 ( .A(\u_div/PartRem[31][4] ), .B(\u_div/u_add_PartRem_2_30/n3 ), 
        .CO(\u_div/u_add_PartRem_2_30/n2 ), .S(\u_div/SumTmp[30][4] ) );
  OR2X1 U99 ( .A(\u_div/PartRem[31][2] ), .B(\u_div/PartRem[31][3] ), .Y(
        \u_div/u_add_PartRem_2_30/n3 ) );
  ADDHXL U100 ( .A(\u_div/PartRem[33][4] ), .B(\u_div/u_add_PartRem_2_32/n3 ), 
        .CO(\u_div/u_add_PartRem_2_32/n2 ), .S(\u_div/SumTmp[32][4] ) );
  ADDHXL U101 ( .A(\u_div/PartRem[32][4] ), .B(\u_div/u_add_PartRem_2_31/n3 ), 
        .CO(\u_div/u_add_PartRem_2_31/n2 ), .S(\u_div/SumTmp[31][4] ) );
  OR2X1 U102 ( .A(\u_div/PartRem[32][2] ), .B(\u_div/PartRem[32][3] ), .Y(
        \u_div/u_add_PartRem_2_31/n3 ) );
  ADDHXL U103 ( .A(\u_div/PartRem[34][4] ), .B(\u_div/u_add_PartRem_2_33/n3 ), 
        .CO(\u_div/u_add_PartRem_2_33/n2 ), .S(\u_div/SumTmp[33][4] ) );
  OR2X1 U104 ( .A(\u_div/PartRem[34][2] ), .B(\u_div/PartRem[34][3] ), .Y(
        \u_div/u_add_PartRem_2_33/n3 ) );
  ADDHXL U105 ( .A(\u_div/PartRem[35][4] ), .B(\u_div/u_add_PartRem_2_34/n3 ), 
        .CO(\u_div/u_add_PartRem_2_34/n2 ), .S(\u_div/SumTmp[34][4] ) );
  OR2X1 U106 ( .A(\u_div/PartRem[35][2] ), .B(\u_div/PartRem[35][3] ), .Y(
        \u_div/u_add_PartRem_2_34/n3 ) );
  ADDHXL U107 ( .A(\u_div/PartRem[36][4] ), .B(\u_div/u_add_PartRem_2_35/n3 ), 
        .CO(\u_div/u_add_PartRem_2_35/n2 ), .S(\u_div/SumTmp[35][4] ) );
  OR2X1 U108 ( .A(\u_div/PartRem[36][2] ), .B(\u_div/PartRem[36][3] ), .Y(
        \u_div/u_add_PartRem_2_35/n3 ) );
  ADDHXL U109 ( .A(\u_div/PartRem[37][4] ), .B(\u_div/u_add_PartRem_2_36/n3 ), 
        .CO(\u_div/u_add_PartRem_2_36/n2 ), .S(\u_div/SumTmp[36][4] ) );
  OR2X1 U110 ( .A(\u_div/PartRem[37][2] ), .B(\u_div/PartRem[37][3] ), .Y(
        \u_div/u_add_PartRem_2_36/n3 ) );
  ADDHXL U111 ( .A(\u_div/PartRem[38][4] ), .B(\u_div/u_add_PartRem_2_37/n3 ), 
        .CO(\u_div/u_add_PartRem_2_37/n2 ), .S(\u_div/SumTmp[37][4] ) );
  ADDHXL U112 ( .A(\u_div/PartRem[39][4] ), .B(\u_div/u_add_PartRem_2_38/n3 ), 
        .CO(\u_div/u_add_PartRem_2_38/n2 ), .S(\u_div/SumTmp[38][4] ) );
  OR2X1 U113 ( .A(\u_div/PartRem[39][2] ), .B(\u_div/PartRem[39][3] ), .Y(
        \u_div/u_add_PartRem_2_38/n3 ) );
  OR2X1 U114 ( .A(\u_div/PartRem[40][2] ), .B(\u_div/PartRem[40][3] ), .Y(
        \u_div/u_add_PartRem_2_39/n3 ) );
  ADDHXL U115 ( .A(\u_div/PartRem[41][4] ), .B(\u_div/u_add_PartRem_2_40/n3 ), 
        .CO(\u_div/u_add_PartRem_2_40/n2 ), .S(\u_div/SumTmp[40][4] ) );
  OR2X1 U116 ( .A(\u_div/PartRem[41][2] ), .B(\u_div/PartRem[41][3] ), .Y(
        \u_div/u_add_PartRem_2_40/n3 ) );
  ADDHXL U117 ( .A(\u_div/PartRem[42][4] ), .B(\u_div/u_add_PartRem_2_41/n3 ), 
        .CO(\u_div/u_add_PartRem_2_41/n2 ), .S(\u_div/SumTmp[41][4] ) );
  OR2X1 U118 ( .A(\u_div/PartRem[42][2] ), .B(\u_div/PartRem[42][3] ), .Y(
        \u_div/u_add_PartRem_2_41/n3 ) );
  ADDHXL U119 ( .A(\u_div/PartRem[43][4] ), .B(\u_div/u_add_PartRem_2_42/n3 ), 
        .CO(\u_div/u_add_PartRem_2_42/n2 ), .S(\u_div/SumTmp[42][4] ) );
  ADDHXL U120 ( .A(\u_div/PartRem[44][4] ), .B(\u_div/u_add_PartRem_2_43/n3 ), 
        .CO(\u_div/u_add_PartRem_2_43/n2 ), .S(\u_div/SumTmp[43][4] ) );
  OR2X1 U121 ( .A(\u_div/PartRem[44][2] ), .B(\u_div/PartRem[44][3] ), .Y(
        \u_div/u_add_PartRem_2_43/n3 ) );
  ADDHXL U122 ( .A(\u_div/PartRem[45][4] ), .B(\u_div/u_add_PartRem_2_44/n3 ), 
        .CO(\u_div/u_add_PartRem_2_44/n2 ), .S(\u_div/SumTmp[44][4] ) );
  OR2X1 U123 ( .A(\u_div/PartRem[45][2] ), .B(\u_div/PartRem[45][3] ), .Y(
        \u_div/u_add_PartRem_2_44/n3 ) );
  ADDHXL U124 ( .A(\u_div/PartRem[46][4] ), .B(\u_div/u_add_PartRem_2_45/n3 ), 
        .CO(\u_div/u_add_PartRem_2_45/n2 ), .S(\u_div/SumTmp[45][4] ) );
  OR2X1 U125 ( .A(\u_div/PartRem[46][2] ), .B(\u_div/PartRem[46][3] ), .Y(
        \u_div/u_add_PartRem_2_45/n3 ) );
  ADDHXL U126 ( .A(\u_div/PartRem[47][4] ), .B(\u_div/u_add_PartRem_2_46/n3 ), 
        .CO(\u_div/u_add_PartRem_2_46/n2 ), .S(\u_div/SumTmp[46][4] ) );
  OR2X1 U127 ( .A(\u_div/PartRem[47][2] ), .B(\u_div/PartRem[47][3] ), .Y(
        \u_div/u_add_PartRem_2_46/n3 ) );
  ADDHXL U128 ( .A(\u_div/PartRem[48][4] ), .B(\u_div/u_add_PartRem_2_47/n3 ), 
        .CO(\u_div/u_add_PartRem_2_47/n2 ), .S(\u_div/SumTmp[47][4] ) );
  ADDHXL U129 ( .A(\u_div/PartRem[50][4] ), .B(\u_div/u_add_PartRem_2_49/n3 ), 
        .CO(\u_div/u_add_PartRem_2_49/n2 ), .S(\u_div/SumTmp[49][4] ) );
  OR2X1 U130 ( .A(\u_div/PartRem[50][2] ), .B(\u_div/PartRem[50][3] ), .Y(
        \u_div/u_add_PartRem_2_49/n3 ) );
  ADDHXL U131 ( .A(\u_div/PartRem[49][4] ), .B(\u_div/u_add_PartRem_2_48/n3 ), 
        .CO(\u_div/u_add_PartRem_2_48/n2 ), .S(\u_div/SumTmp[48][4] ) );
  OR2X1 U132 ( .A(\u_div/PartRem[49][2] ), .B(\u_div/PartRem[49][3] ), .Y(
        \u_div/u_add_PartRem_2_48/n3 ) );
  ADDHXL U133 ( .A(\u_div/PartRem[51][4] ), .B(\u_div/u_add_PartRem_2_50/n3 ), 
        .CO(\u_div/u_add_PartRem_2_50/n2 ), .S(\u_div/SumTmp[50][4] ) );
  OR2X1 U134 ( .A(\u_div/PartRem[51][2] ), .B(\u_div/PartRem[51][3] ), .Y(
        \u_div/u_add_PartRem_2_50/n3 ) );
  ADDHXL U135 ( .A(\u_div/PartRem[52][4] ), .B(\u_div/u_add_PartRem_2_51/n3 ), 
        .CO(\u_div/u_add_PartRem_2_51/n2 ), .S(\u_div/SumTmp[51][4] ) );
  OR2X1 U136 ( .A(\u_div/PartRem[52][2] ), .B(\u_div/PartRem[52][3] ), .Y(
        \u_div/u_add_PartRem_2_51/n3 ) );
  ADDHXL U137 ( .A(\u_div/PartRem[53][4] ), .B(\u_div/u_add_PartRem_2_52/n3 ), 
        .CO(\u_div/u_add_PartRem_2_52/n2 ), .S(\u_div/SumTmp[52][4] ) );
  ADDHXL U138 ( .A(\u_div/PartRem[54][4] ), .B(\u_div/u_add_PartRem_2_53/n3 ), 
        .CO(\u_div/u_add_PartRem_2_53/n2 ), .S(\u_div/SumTmp[53][4] ) );
  OR2X1 U139 ( .A(\u_div/PartRem[54][2] ), .B(\u_div/PartRem[54][3] ), .Y(
        \u_div/u_add_PartRem_2_53/n3 ) );
  ADDHXL U140 ( .A(\u_div/PartRem[55][4] ), .B(\u_div/u_add_PartRem_2_54/n3 ), 
        .CO(\u_div/u_add_PartRem_2_54/n2 ), .S(\u_div/SumTmp[54][4] ) );
  OR2X1 U141 ( .A(\u_div/PartRem[55][2] ), .B(\u_div/PartRem[55][3] ), .Y(
        \u_div/u_add_PartRem_2_54/n3 ) );
  ADDHXL U142 ( .A(\u_div/PartRem[56][4] ), .B(\u_div/u_add_PartRem_2_55/n3 ), 
        .CO(\u_div/u_add_PartRem_2_55/n2 ), .S(\u_div/SumTmp[55][4] ) );
  OR2X1 U143 ( .A(\u_div/PartRem[56][2] ), .B(\u_div/PartRem[56][3] ), .Y(
        \u_div/u_add_PartRem_2_55/n3 ) );
  ADDHXL U144 ( .A(\u_div/PartRem[57][4] ), .B(\u_div/u_add_PartRem_2_56/n3 ), 
        .CO(\u_div/u_add_PartRem_2_56/n2 ), .S(\u_div/SumTmp[56][4] ) );
  OR2X1 U145 ( .A(\u_div/PartRem[57][2] ), .B(\u_div/PartRem[57][3] ), .Y(
        \u_div/u_add_PartRem_2_56/n3 ) );
  ADDHXL U146 ( .A(\u_div/PartRem[58][4] ), .B(\u_div/u_add_PartRem_2_57/n3 ), 
        .CO(\u_div/u_add_PartRem_2_57/n2 ), .S(\u_div/SumTmp[57][4] ) );
  OR2X1 U147 ( .A(\u_div/PartRem[58][2] ), .B(\u_div/PartRem[58][3] ), .Y(
        \u_div/u_add_PartRem_2_57/n3 ) );
  NOR2X1 U148 ( .A(\u_div/PartRem[63][0] ), .B(\u_div/PartRem[62][0] ), .Y(n8)
         );
  OR2X1 U149 ( .A(\u_div/PartRem[16][5] ), .B(\u_div/u_add_PartRem_2_15/n2 ), 
        .Y(\u_div/CryTmp[15][6] ) );
  OR2X1 U150 ( .A(\u_div/PartRem[21][5] ), .B(\u_div/u_add_PartRem_2_20/n2 ), 
        .Y(\u_div/CryTmp[20][6] ) );
  ADDHXL U151 ( .A(\u_div/PartRem[2][4] ), .B(\u_div/u_add_PartRem_2_1/n3 ), 
        .CO(\u_div/u_add_PartRem_2_1/n2 ), .S(\u_div/SumTmp[1][4] ) );
  OR2X1 U152 ( .A(\u_div/PartRem[2][2] ), .B(\u_div/PartRem[2][3] ), .Y(
        \u_div/u_add_PartRem_2_1/n3 ) );
  OR2X1 U153 ( .A(\u_div/PartRem[26][5] ), .B(\u_div/u_add_PartRem_2_25/n2 ), 
        .Y(\u_div/CryTmp[25][6] ) );
  OR2X1 U154 ( .A(\u_div/PartRem[31][5] ), .B(\u_div/u_add_PartRem_2_30/n2 ), 
        .Y(\u_div/CryTmp[30][6] ) );
  OR2X1 U155 ( .A(\u_div/PartRem[36][5] ), .B(\u_div/u_add_PartRem_2_35/n2 ), 
        .Y(\u_div/CryTmp[35][6] ) );
  OR2X1 U156 ( .A(\u_div/PartRem[41][5] ), .B(\u_div/u_add_PartRem_2_40/n2 ), 
        .Y(\u_div/CryTmp[40][6] ) );
  OR2X1 U157 ( .A(\u_div/PartRem[46][5] ), .B(\u_div/u_add_PartRem_2_45/n2 ), 
        .Y(\u_div/CryTmp[45][6] ) );
  OR2X1 U158 ( .A(\u_div/PartRem[51][5] ), .B(\u_div/u_add_PartRem_2_50/n2 ), 
        .Y(\u_div/CryTmp[50][6] ) );
  OR2X1 U159 ( .A(\u_div/PartRem[56][5] ), .B(\u_div/u_add_PartRem_2_55/n2 ), 
        .Y(\u_div/CryTmp[55][6] ) );
  NOR2BX2 U160 ( .AN(\u_div/PartRem[64][0] ), .B(n8), .Y(\u_div/CryTmp[59][6] ) );
  AO21X1 U161 ( .A0(\u_div/PartRem[1][4] ), .A1(n6), .B0(\u_div/PartRem[1][5] ), .Y(\u_div/CryTmp[0][6] ) );
  OR2XL U162 ( .A(\u_div/PartRem[59][2] ), .B(\u_div/PartRem[59][3] ), .Y(
        \u_div/u_add_PartRem_2_58/n3 ) );
  XNOR2XL U163 ( .A(\u_div/PartRem[64][0] ), .B(n8), .Y(\u_div/SumTmp[59][4] )
         );
  XOR2XL U164 ( .A(\u_div/CryTmp[59][6] ), .B(n3), .Y(\u_div/QInv[59] ) );
  XOR2XL U165 ( .A(\u_div/CryTmp[1][6] ), .B(n4), .Y(\u_div/QInv[1] ) );
  XOR2XL U166 ( .A(\u_div/CryTmp[54][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[54] ) );
  XOR2XL U167 ( .A(\u_div/CryTmp[55][6] ), .B(n4), .Y(\u_div/QInv[55] ) );
  XOR2XL U168 ( .A(\u_div/CryTmp[51][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[51] ) );
  XOR2XL U169 ( .A(\u_div/CryTmp[52][6] ), .B(n4), .Y(\u_div/QInv[52] ) );
  XOR2XL U170 ( .A(\u_div/CryTmp[47][6] ), .B(n4), .Y(\u_div/QInv[47] ) );
  XOR2XL U171 ( .A(\u_div/CryTmp[44][6] ), .B(n4), .Y(\u_div/QInv[44] ) );
  XOR2XL U172 ( .A(\u_div/CryTmp[41][6] ), .B(n4), .Y(\u_div/QInv[41] ) );
  XOR2XL U173 ( .A(\u_div/CryTmp[34][6] ), .B(n4), .Y(\u_div/QInv[34] ) );
  XOR2XL U174 ( .A(\u_div/CryTmp[36][6] ), .B(n4), .Y(\u_div/QInv[36] ) );
  XOR2XL U175 ( .A(\u_div/CryTmp[31][6] ), .B(n4), .Y(\u_div/QInv[31] ) );
  XOR2XL U176 ( .A(\u_div/CryTmp[26][6] ), .B(n4), .Y(\u_div/QInv[26] ) );
  XOR2XL U177 ( .A(\u_div/CryTmp[22][6] ), .B(n5), .Y(\u_div/QInv[22] ) );
  XOR2XL U178 ( .A(\u_div/CryTmp[23][6] ), .B(n4), .Y(\u_div/QInv[23] ) );
  XOR2XL U179 ( .A(\u_div/CryTmp[20][6] ), .B(n4), .Y(\u_div/QInv[20] ) );
  XOR2XL U180 ( .A(\u_div/CryTmp[14][6] ), .B(n4), .Y(\u_div/QInv[14] ) );
  XOR2XL U181 ( .A(\u_div/CryTmp[12][6] ), .B(n4), .Y(\u_div/QInv[12] ) );
  XOR2XL U182 ( .A(\u_div/CryTmp[11][6] ), .B(n4), .Y(\u_div/QInv[11] ) );
  XOR2XL U183 ( .A(\u_div/CryTmp[4][6] ), .B(n4), .Y(\u_div/QInv[4] ) );
  XOR2XL U184 ( .A(\u_div/CryTmp[57][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[57] ) );
  XOR2XL U185 ( .A(\u_div/CryTmp[50][6] ), .B(n3), .Y(\u_div/QInv[50] ) );
  XOR2XL U186 ( .A(\u_div/CryTmp[45][6] ), .B(n3), .Y(\u_div/QInv[45] ) );
  XOR2XL U187 ( .A(\u_div/CryTmp[46][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[46] ) );
  XOR2XL U188 ( .A(\u_div/CryTmp[42][6] ), .B(n3), .Y(\u_div/QInv[42] ) );
  XOR2XL U189 ( .A(\u_div/CryTmp[43][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[43] ) );
  XOR2XL U190 ( .A(\u_div/CryTmp[40][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[40] ) );
  XOR2XL U191 ( .A(\u_div/CryTmp[37][6] ), .B(n3), .Y(\u_div/QInv[37] ) );
  XOR2XL U192 ( .A(\u_div/CryTmp[35][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[35] ) );
  XOR2XL U193 ( .A(\u_div/CryTmp[33][6] ), .B(n5), .Y(\u_div/QInv[33] ) );
  XOR2XL U194 ( .A(\u_div/CryTmp[32][6] ), .B(n3), .Y(\u_div/QInv[32] ) );
  XOR2XL U195 ( .A(\u_div/CryTmp[30][6] ), .B(n5), .Y(\u_div/QInv[30] ) );
  XOR2XL U196 ( .A(\u_div/CryTmp[27][6] ), .B(n3), .Y(\u_div/QInv[27] ) );
  XOR2XL U197 ( .A(\u_div/CryTmp[25][6] ), .B(n5), .Y(\u_div/QInv[25] ) );
  XOR2XL U198 ( .A(\u_div/CryTmp[24][6] ), .B(n3), .Y(\u_div/QInv[24] ) );
  XOR2XL U199 ( .A(\u_div/CryTmp[21][6] ), .B(n3), .Y(\u_div/QInv[21] ) );
  XOR2XL U200 ( .A(\u_div/CryTmp[17][6] ), .B(n5), .Y(\u_div/QInv[17] ) );
  XOR2XL U201 ( .A(\u_div/CryTmp[16][6] ), .B(n4), .Y(\u_div/QInv[16] ) );
  XOR2XL U202 ( .A(\u_div/CryTmp[15][6] ), .B(n3), .Y(\u_div/QInv[15] ) );
  XOR2XL U203 ( .A(\u_div/CryTmp[13][6] ), .B(n4), .Y(\u_div/QInv[13] ) );
  XOR2XL U204 ( .A(\u_div/CryTmp[5][6] ), .B(n4), .Y(\u_div/QInv[5] ) );
  XOR2XL U205 ( .A(\u_div/CryTmp[6][6] ), .B(n4), .Y(\u_div/QInv[6] ) );
  XOR2XL U206 ( .A(\u_div/CryTmp[7][6] ), .B(n4), .Y(\u_div/QInv[7] ) );
  XOR2XL U207 ( .A(\u_div/CryTmp[10][6] ), .B(n4), .Y(\u_div/QInv[10] ) );
  XOR2XL U208 ( .A(\u_div/CryTmp[2][6] ), .B(n3), .Y(\u_div/QInv[2] ) );
  XOR2XL U209 ( .A(\u_div/CryTmp[3][6] ), .B(n3), .Y(\u_div/QInv[3] ) );
  INVXL U210 ( .A(\u_div/PartRem[59][2] ), .Y(\u_div/SumTmp[58][2] ) );
  INVXL U211 ( .A(\u_div/PartRem[55][2] ), .Y(\u_div/SumTmp[54][2] ) );
  INVXL U212 ( .A(\u_div/PartRem[50][2] ), .Y(\u_div/SumTmp[49][2] ) );
  INVXL U213 ( .A(\u_div/PartRem[45][2] ), .Y(\u_div/SumTmp[44][2] ) );
  INVXL U214 ( .A(\u_div/PartRem[40][2] ), .Y(\u_div/SumTmp[39][2] ) );
  INVXL U215 ( .A(\u_div/PartRem[35][2] ), .Y(\u_div/SumTmp[34][2] ) );
  INVXL U216 ( .A(\u_div/PartRem[30][2] ), .Y(\u_div/SumTmp[29][2] ) );
  INVXL U217 ( .A(\u_div/PartRem[25][2] ), .Y(\u_div/SumTmp[24][2] ) );
  INVXL U218 ( .A(\u_div/PartRem[20][2] ), .Y(\u_div/SumTmp[19][2] ) );
  INVXL U219 ( .A(\u_div/PartRem[15][2] ), .Y(\u_div/SumTmp[14][2] ) );
  INVXL U220 ( .A(\u_div/PartRem[10][2] ), .Y(\u_div/SumTmp[9][2] ) );
  INVXL U221 ( .A(\u_div/PartRem[5][2] ), .Y(\u_div/SumTmp[4][2] ) );
  INVX3 U222 ( .A(n2), .Y(n3) );
  MXI2X1 U223 ( .A(\u_div/SumTmp[1][1] ), .B(\u_div/SumTmp[1][1] ), .S0(
        \u_div/CryTmp[1][6] ), .Y(n1) );
  CLKINVX1 U224 ( .A(n5), .Y(n2) );
  MXI2X1 U225 ( .A(n7), .B(\u_div/PartRem[62][0] ), .S0(\u_div/CryTmp[59][6] ), 
        .Y(\u_div/PartRem[59][3] ) );
  CLKINVX1 U226 ( .A(\u_div/PartRem[62][0] ), .Y(n7) );
  MXI2X1 U227 ( .A(\u_div/SumTmp[58][2] ), .B(\u_div/PartRem[59][2] ), .S0(
        \u_div/CryTmp[58][6] ), .Y(\u_div/PartRem[58][3] ) );
  MXI2X1 U228 ( .A(\u_div/SumTmp[57][2] ), .B(\u_div/PartRem[58][2] ), .S0(
        \u_div/CryTmp[57][6] ), .Y(\u_div/PartRem[57][3] ) );
  CLKINVX1 U229 ( .A(\u_div/PartRem[58][2] ), .Y(\u_div/SumTmp[57][2] ) );
  CLKINVX1 U230 ( .A(\u_div/PartRem[57][2] ), .Y(\u_div/SumTmp[56][2] ) );
  MXI2X1 U231 ( .A(\u_div/SumTmp[54][2] ), .B(\u_div/PartRem[55][2] ), .S0(
        \u_div/CryTmp[54][6] ), .Y(\u_div/PartRem[54][3] ) );
  CLKINVX1 U232 ( .A(\u_div/PartRem[54][2] ), .Y(\u_div/SumTmp[53][2] ) );
  MXI2X1 U233 ( .A(\u_div/SumTmp[52][2] ), .B(\u_div/PartRem[53][2] ), .S0(
        \u_div/CryTmp[52][6] ), .Y(\u_div/PartRem[52][3] ) );
  CLKINVX1 U234 ( .A(\u_div/PartRem[53][2] ), .Y(\u_div/SumTmp[52][2] ) );
  MXI2X1 U235 ( .A(\u_div/SumTmp[51][2] ), .B(\u_div/PartRem[52][2] ), .S0(
        \u_div/CryTmp[51][6] ), .Y(\u_div/PartRem[51][3] ) );
  CLKINVX1 U236 ( .A(\u_div/PartRem[52][2] ), .Y(\u_div/SumTmp[51][2] ) );
  CLKINVX1 U237 ( .A(\u_div/PartRem[49][2] ), .Y(\u_div/SumTmp[48][2] ) );
  MXI2X1 U238 ( .A(\u_div/SumTmp[47][2] ), .B(\u_div/PartRem[48][2] ), .S0(
        \u_div/CryTmp[47][6] ), .Y(\u_div/PartRem[47][3] ) );
  CLKINVX1 U239 ( .A(\u_div/PartRem[48][2] ), .Y(\u_div/SumTmp[47][2] ) );
  MXI2X1 U240 ( .A(\u_div/SumTmp[46][2] ), .B(\u_div/PartRem[47][2] ), .S0(
        \u_div/CryTmp[46][6] ), .Y(\u_div/PartRem[46][3] ) );
  CLKINVX1 U241 ( .A(\u_div/PartRem[47][2] ), .Y(\u_div/SumTmp[46][2] ) );
  MXI2X1 U242 ( .A(\u_div/SumTmp[44][2] ), .B(\u_div/PartRem[45][2] ), .S0(
        \u_div/CryTmp[44][6] ), .Y(\u_div/PartRem[44][3] ) );
  CLKINVX1 U243 ( .A(\u_div/PartRem[44][2] ), .Y(\u_div/SumTmp[43][2] ) );
  MXI2X1 U244 ( .A(\u_div/SumTmp[42][2] ), .B(\u_div/PartRem[43][2] ), .S0(
        \u_div/CryTmp[42][6] ), .Y(\u_div/PartRem[42][3] ) );
  CLKINVX1 U245 ( .A(\u_div/PartRem[43][2] ), .Y(\u_div/SumTmp[42][2] ) );
  MXI2X1 U246 ( .A(\u_div/SumTmp[41][2] ), .B(\u_div/PartRem[42][2] ), .S0(
        \u_div/CryTmp[41][6] ), .Y(\u_div/PartRem[41][3] ) );
  CLKINVX1 U247 ( .A(\u_div/PartRem[42][2] ), .Y(\u_div/SumTmp[41][2] ) );
  MXI2X1 U248 ( .A(\u_div/SumTmp[39][2] ), .B(\u_div/PartRem[40][2] ), .S0(
        \u_div/CryTmp[39][6] ), .Y(\u_div/PartRem[39][3] ) );
  CLKINVX1 U249 ( .A(\u_div/PartRem[39][2] ), .Y(\u_div/SumTmp[38][2] ) );
  MXI2X1 U250 ( .A(\u_div/SumTmp[37][2] ), .B(\u_div/PartRem[38][2] ), .S0(
        \u_div/CryTmp[37][6] ), .Y(\u_div/PartRem[37][3] ) );
  CLKINVX1 U251 ( .A(\u_div/PartRem[38][2] ), .Y(\u_div/SumTmp[37][2] ) );
  MXI2X1 U252 ( .A(\u_div/SumTmp[36][2] ), .B(\u_div/PartRem[37][2] ), .S0(
        \u_div/CryTmp[36][6] ), .Y(\u_div/PartRem[36][3] ) );
  CLKINVX1 U253 ( .A(\u_div/PartRem[37][2] ), .Y(\u_div/SumTmp[36][2] ) );
  MXI2X1 U254 ( .A(\u_div/SumTmp[34][2] ), .B(\u_div/PartRem[35][2] ), .S0(
        \u_div/CryTmp[34][6] ), .Y(\u_div/PartRem[34][3] ) );
  CLKINVX1 U255 ( .A(\u_div/PartRem[34][2] ), .Y(\u_div/SumTmp[33][2] ) );
  MXI2X1 U256 ( .A(\u_div/SumTmp[32][2] ), .B(\u_div/PartRem[33][2] ), .S0(
        \u_div/CryTmp[32][6] ), .Y(\u_div/PartRem[32][3] ) );
  CLKINVX1 U257 ( .A(\u_div/PartRem[33][2] ), .Y(\u_div/SumTmp[32][2] ) );
  MXI2X1 U258 ( .A(\u_div/SumTmp[31][2] ), .B(\u_div/PartRem[32][2] ), .S0(
        \u_div/CryTmp[31][6] ), .Y(\u_div/PartRem[31][3] ) );
  CLKINVX1 U259 ( .A(\u_div/PartRem[32][2] ), .Y(\u_div/SumTmp[31][2] ) );
  MXI2X1 U260 ( .A(\u_div/SumTmp[29][2] ), .B(\u_div/PartRem[30][2] ), .S0(
        \u_div/CryTmp[29][6] ), .Y(\u_div/PartRem[29][3] ) );
  CLKINVX1 U261 ( .A(\u_div/PartRem[29][2] ), .Y(\u_div/SumTmp[28][2] ) );
  MXI2X1 U262 ( .A(\u_div/SumTmp[27][2] ), .B(\u_div/PartRem[28][2] ), .S0(
        \u_div/CryTmp[27][6] ), .Y(\u_div/PartRem[27][3] ) );
  CLKINVX1 U263 ( .A(\u_div/PartRem[28][2] ), .Y(\u_div/SumTmp[27][2] ) );
  MXI2X1 U264 ( .A(\u_div/SumTmp[26][2] ), .B(\u_div/PartRem[27][2] ), .S0(
        \u_div/CryTmp[26][6] ), .Y(\u_div/PartRem[26][3] ) );
  CLKINVX1 U265 ( .A(\u_div/PartRem[27][2] ), .Y(\u_div/SumTmp[26][2] ) );
  MXI2X1 U266 ( .A(\u_div/SumTmp[24][2] ), .B(\u_div/PartRem[25][2] ), .S0(
        \u_div/CryTmp[24][6] ), .Y(\u_div/PartRem[24][3] ) );
  CLKINVX1 U267 ( .A(\u_div/PartRem[24][2] ), .Y(\u_div/SumTmp[23][2] ) );
  MXI2X1 U268 ( .A(\u_div/SumTmp[22][2] ), .B(\u_div/PartRem[23][2] ), .S0(
        \u_div/CryTmp[22][6] ), .Y(\u_div/PartRem[22][3] ) );
  CLKINVX1 U269 ( .A(\u_div/PartRem[23][2] ), .Y(\u_div/SumTmp[22][2] ) );
  MXI2X1 U270 ( .A(\u_div/SumTmp[21][2] ), .B(\u_div/PartRem[22][2] ), .S0(
        \u_div/CryTmp[21][6] ), .Y(\u_div/PartRem[21][3] ) );
  CLKINVX1 U271 ( .A(\u_div/PartRem[22][2] ), .Y(\u_div/SumTmp[21][2] ) );
  CLKINVX1 U272 ( .A(\u_div/PartRem[19][2] ), .Y(\u_div/SumTmp[18][2] ) );
  MXI2X1 U273 ( .A(\u_div/SumTmp[17][2] ), .B(\u_div/PartRem[18][2] ), .S0(
        \u_div/CryTmp[17][6] ), .Y(\u_div/PartRem[17][3] ) );
  CLKINVX1 U274 ( .A(\u_div/PartRem[18][2] ), .Y(\u_div/SumTmp[17][2] ) );
  MXI2X1 U275 ( .A(\u_div/SumTmp[16][2] ), .B(\u_div/PartRem[17][2] ), .S0(
        \u_div/CryTmp[16][6] ), .Y(\u_div/PartRem[16][3] ) );
  CLKINVX1 U276 ( .A(\u_div/PartRem[17][2] ), .Y(\u_div/SumTmp[16][2] ) );
  MXI2X1 U277 ( .A(\u_div/SumTmp[14][2] ), .B(\u_div/PartRem[15][2] ), .S0(
        \u_div/CryTmp[14][6] ), .Y(\u_div/PartRem[14][3] ) );
  CLKINVX1 U278 ( .A(\u_div/PartRem[14][2] ), .Y(\u_div/SumTmp[13][2] ) );
  MXI2X1 U279 ( .A(\u_div/SumTmp[12][2] ), .B(\u_div/PartRem[13][2] ), .S0(
        \u_div/CryTmp[12][6] ), .Y(\u_div/PartRem[12][3] ) );
  CLKINVX1 U280 ( .A(\u_div/PartRem[13][2] ), .Y(\u_div/SumTmp[12][2] ) );
  MXI2X1 U281 ( .A(\u_div/SumTmp[11][2] ), .B(\u_div/PartRem[12][2] ), .S0(
        \u_div/CryTmp[11][6] ), .Y(\u_div/PartRem[11][3] ) );
  CLKINVX1 U282 ( .A(\u_div/PartRem[12][2] ), .Y(\u_div/SumTmp[11][2] ) );
  CLKINVX1 U283 ( .A(\u_div/PartRem[9][2] ), .Y(\u_div/SumTmp[8][2] ) );
  CLKINVX1 U284 ( .A(\u_div/PartRem[8][2] ), .Y(\u_div/SumTmp[7][2] ) );
  MXI2X1 U285 ( .A(\u_div/SumTmp[6][2] ), .B(\u_div/PartRem[7][2] ), .S0(
        \u_div/CryTmp[6][6] ), .Y(\u_div/PartRem[6][3] ) );
  CLKINVX1 U286 ( .A(\u_div/PartRem[7][2] ), .Y(\u_div/SumTmp[6][2] ) );
  MXI2X1 U287 ( .A(\u_div/SumTmp[4][2] ), .B(\u_div/PartRem[5][2] ), .S0(
        \u_div/CryTmp[4][6] ), .Y(\u_div/PartRem[4][3] ) );
  CLKINVX1 U288 ( .A(\u_div/PartRem[4][2] ), .Y(\u_div/SumTmp[3][2] ) );
  MXI2X1 U289 ( .A(\u_div/SumTmp[2][2] ), .B(\u_div/PartRem[3][2] ), .S0(
        \u_div/CryTmp[2][6] ), .Y(\u_div/PartRem[2][3] ) );
  CLKINVX1 U290 ( .A(\u_div/PartRem[3][2] ), .Y(\u_div/SumTmp[2][2] ) );
  MXI2X1 U291 ( .A(\u_div/SumTmp[55][2] ), .B(\u_div/PartRem[56][2] ), .S0(
        \u_div/CryTmp[55][6] ), .Y(\u_div/PartRem[55][3] ) );
  CLKINVX1 U292 ( .A(\u_div/PartRem[56][2] ), .Y(\u_div/SumTmp[55][2] ) );
  MXI2X1 U293 ( .A(\u_div/SumTmp[50][2] ), .B(\u_div/PartRem[51][2] ), .S0(
        \u_div/CryTmp[50][6] ), .Y(\u_div/PartRem[50][3] ) );
  CLKINVX1 U294 ( .A(\u_div/PartRem[51][2] ), .Y(\u_div/SumTmp[50][2] ) );
  MXI2X1 U295 ( .A(\u_div/SumTmp[45][2] ), .B(\u_div/PartRem[46][2] ), .S0(
        \u_div/CryTmp[45][6] ), .Y(\u_div/PartRem[45][3] ) );
  CLKINVX1 U296 ( .A(\u_div/PartRem[46][2] ), .Y(\u_div/SumTmp[45][2] ) );
  MXI2X1 U297 ( .A(\u_div/SumTmp[40][2] ), .B(\u_div/PartRem[41][2] ), .S0(
        \u_div/CryTmp[40][6] ), .Y(\u_div/PartRem[40][3] ) );
  CLKINVX1 U298 ( .A(\u_div/PartRem[41][2] ), .Y(\u_div/SumTmp[40][2] ) );
  MXI2X1 U299 ( .A(\u_div/SumTmp[35][2] ), .B(\u_div/PartRem[36][2] ), .S0(
        \u_div/CryTmp[35][6] ), .Y(\u_div/PartRem[35][3] ) );
  CLKINVX1 U300 ( .A(\u_div/PartRem[36][2] ), .Y(\u_div/SumTmp[35][2] ) );
  MXI2X1 U301 ( .A(\u_div/SumTmp[30][2] ), .B(\u_div/PartRem[31][2] ), .S0(
        \u_div/CryTmp[30][6] ), .Y(\u_div/PartRem[30][3] ) );
  CLKINVX1 U302 ( .A(\u_div/PartRem[31][2] ), .Y(\u_div/SumTmp[30][2] ) );
  MXI2X1 U303 ( .A(\u_div/SumTmp[25][2] ), .B(\u_div/PartRem[26][2] ), .S0(
        \u_div/CryTmp[25][6] ), .Y(\u_div/PartRem[25][3] ) );
  CLKINVX1 U304 ( .A(\u_div/PartRem[26][2] ), .Y(\u_div/SumTmp[25][2] ) );
  MXI2X1 U305 ( .A(\u_div/SumTmp[20][2] ), .B(\u_div/PartRem[21][2] ), .S0(
        \u_div/CryTmp[20][6] ), .Y(\u_div/PartRem[20][3] ) );
  CLKINVX1 U306 ( .A(\u_div/PartRem[21][2] ), .Y(\u_div/SumTmp[20][2] ) );
  MXI2X1 U307 ( .A(\u_div/SumTmp[15][2] ), .B(\u_div/PartRem[16][2] ), .S0(
        \u_div/CryTmp[15][6] ), .Y(\u_div/PartRem[15][3] ) );
  CLKINVX1 U308 ( .A(\u_div/PartRem[16][2] ), .Y(\u_div/SumTmp[15][2] ) );
  MXI2X1 U309 ( .A(\u_div/SumTmp[10][2] ), .B(\u_div/PartRem[11][2] ), .S0(
        \u_div/CryTmp[10][6] ), .Y(\u_div/PartRem[10][3] ) );
  CLKINVX1 U310 ( .A(\u_div/PartRem[11][2] ), .Y(\u_div/SumTmp[10][2] ) );
  MXI2X1 U311 ( .A(\u_div/SumTmp[5][2] ), .B(\u_div/PartRem[6][2] ), .S0(
        \u_div/CryTmp[5][6] ), .Y(\u_div/PartRem[5][3] ) );
  CLKINVX1 U312 ( .A(\u_div/PartRem[6][2] ), .Y(\u_div/SumTmp[5][2] ) );
  CLKINVX1 U313 ( .A(\u_div/PartRem[2][2] ), .Y(\u_div/SumTmp[1][2] ) );
  INVX4 U314 ( .A(n2), .Y(n4) );
  CLKBUFX3 U315 ( .A(\u_div/QInv[63] ), .Y(n5) );
  XNOR2X1 U316 ( .A(\u_div/PartRem[59][3] ), .B(\u_div/PartRem[59][2] ), .Y(
        \u_div/SumTmp[58][3] ) );
  OR2X1 U317 ( .A(\u_div/PartRem[58][5] ), .B(\u_div/u_add_PartRem_2_57/n2 ), 
        .Y(\u_div/CryTmp[57][6] ) );
  XNOR2X1 U318 ( .A(\u_div/PartRem[58][3] ), .B(\u_div/PartRem[58][2] ), .Y(
        \u_div/SumTmp[57][3] ) );
  XNOR2X1 U319 ( .A(\u_div/PartRem[57][3] ), .B(\u_div/PartRem[57][2] ), .Y(
        \u_div/SumTmp[56][3] ) );
  XNOR2X1 U320 ( .A(\u_div/PartRem[56][3] ), .B(\u_div/PartRem[56][2] ), .Y(
        \u_div/SumTmp[55][3] ) );
  OR2X1 U321 ( .A(\u_div/PartRem[55][5] ), .B(\u_div/u_add_PartRem_2_54/n2 ), 
        .Y(\u_div/CryTmp[54][6] ) );
  XNOR2X1 U322 ( .A(\u_div/PartRem[55][3] ), .B(\u_div/PartRem[55][2] ), .Y(
        \u_div/SumTmp[54][3] ) );
  XNOR2X1 U323 ( .A(\u_div/PartRem[54][3] ), .B(\u_div/PartRem[54][2] ), .Y(
        \u_div/SumTmp[53][3] ) );
  OR2X1 U324 ( .A(\u_div/PartRem[53][5] ), .B(\u_div/u_add_PartRem_2_52/n2 ), 
        .Y(\u_div/CryTmp[52][6] ) );
  XNOR2X1 U325 ( .A(\u_div/PartRem[53][3] ), .B(\u_div/PartRem[53][2] ), .Y(
        \u_div/SumTmp[52][3] ) );
  OR2X1 U326 ( .A(\u_div/PartRem[53][2] ), .B(\u_div/PartRem[53][3] ), .Y(
        \u_div/u_add_PartRem_2_52/n3 ) );
  OR2X1 U327 ( .A(\u_div/PartRem[52][5] ), .B(\u_div/u_add_PartRem_2_51/n2 ), 
        .Y(\u_div/CryTmp[51][6] ) );
  XNOR2X1 U328 ( .A(\u_div/PartRem[52][3] ), .B(\u_div/PartRem[52][2] ), .Y(
        \u_div/SumTmp[51][3] ) );
  XNOR2X1 U329 ( .A(\u_div/PartRem[51][3] ), .B(\u_div/PartRem[51][2] ), .Y(
        \u_div/SumTmp[50][3] ) );
  XNOR2X1 U330 ( .A(\u_div/PartRem[50][3] ), .B(\u_div/PartRem[50][2] ), .Y(
        \u_div/SumTmp[49][3] ) );
  XNOR2X1 U331 ( .A(\u_div/PartRem[49][3] ), .B(\u_div/PartRem[49][2] ), .Y(
        \u_div/SumTmp[48][3] ) );
  OR2X1 U332 ( .A(\u_div/PartRem[48][5] ), .B(\u_div/u_add_PartRem_2_47/n2 ), 
        .Y(\u_div/CryTmp[47][6] ) );
  XNOR2X1 U333 ( .A(\u_div/PartRem[48][3] ), .B(\u_div/PartRem[48][2] ), .Y(
        \u_div/SumTmp[47][3] ) );
  OR2X1 U334 ( .A(\u_div/PartRem[48][2] ), .B(\u_div/PartRem[48][3] ), .Y(
        \u_div/u_add_PartRem_2_47/n3 ) );
  OR2X1 U335 ( .A(\u_div/PartRem[47][5] ), .B(\u_div/u_add_PartRem_2_46/n2 ), 
        .Y(\u_div/CryTmp[46][6] ) );
  XNOR2X1 U336 ( .A(\u_div/PartRem[47][3] ), .B(\u_div/PartRem[47][2] ), .Y(
        \u_div/SumTmp[46][3] ) );
  XNOR2X1 U337 ( .A(\u_div/PartRem[46][3] ), .B(\u_div/PartRem[46][2] ), .Y(
        \u_div/SumTmp[45][3] ) );
  OR2X1 U338 ( .A(\u_div/PartRem[45][5] ), .B(\u_div/u_add_PartRem_2_44/n2 ), 
        .Y(\u_div/CryTmp[44][6] ) );
  XNOR2X1 U339 ( .A(\u_div/PartRem[45][3] ), .B(\u_div/PartRem[45][2] ), .Y(
        \u_div/SumTmp[44][3] ) );
  OR2X1 U340 ( .A(\u_div/PartRem[44][5] ), .B(\u_div/u_add_PartRem_2_43/n2 ), 
        .Y(\u_div/CryTmp[43][6] ) );
  XNOR2X1 U341 ( .A(\u_div/PartRem[44][3] ), .B(\u_div/PartRem[44][2] ), .Y(
        \u_div/SumTmp[43][3] ) );
  OR2X1 U342 ( .A(\u_div/PartRem[43][5] ), .B(\u_div/u_add_PartRem_2_42/n2 ), 
        .Y(\u_div/CryTmp[42][6] ) );
  XNOR2X1 U343 ( .A(\u_div/PartRem[43][3] ), .B(\u_div/PartRem[43][2] ), .Y(
        \u_div/SumTmp[42][3] ) );
  OR2X1 U344 ( .A(\u_div/PartRem[43][2] ), .B(\u_div/PartRem[43][3] ), .Y(
        \u_div/u_add_PartRem_2_42/n3 ) );
  OR2X1 U345 ( .A(\u_div/PartRem[42][5] ), .B(\u_div/u_add_PartRem_2_41/n2 ), 
        .Y(\u_div/CryTmp[41][6] ) );
  XNOR2X1 U346 ( .A(\u_div/PartRem[42][3] ), .B(\u_div/PartRem[42][2] ), .Y(
        \u_div/SumTmp[41][3] ) );
  XNOR2X1 U347 ( .A(\u_div/PartRem[41][3] ), .B(\u_div/PartRem[41][2] ), .Y(
        \u_div/SumTmp[40][3] ) );
  XNOR2X1 U348 ( .A(\u_div/PartRem[40][3] ), .B(\u_div/PartRem[40][2] ), .Y(
        \u_div/SumTmp[39][3] ) );
  XNOR2X1 U349 ( .A(\u_div/PartRem[39][3] ), .B(\u_div/PartRem[39][2] ), .Y(
        \u_div/SumTmp[38][3] ) );
  OR2X1 U350 ( .A(\u_div/PartRem[38][5] ), .B(\u_div/u_add_PartRem_2_37/n2 ), 
        .Y(\u_div/CryTmp[37][6] ) );
  XNOR2X1 U351 ( .A(\u_div/PartRem[38][3] ), .B(\u_div/PartRem[38][2] ), .Y(
        \u_div/SumTmp[37][3] ) );
  OR2X1 U352 ( .A(\u_div/PartRem[38][2] ), .B(\u_div/PartRem[38][3] ), .Y(
        \u_div/u_add_PartRem_2_37/n3 ) );
  OR2X1 U353 ( .A(\u_div/PartRem[37][5] ), .B(\u_div/u_add_PartRem_2_36/n2 ), 
        .Y(\u_div/CryTmp[36][6] ) );
  XNOR2X1 U354 ( .A(\u_div/PartRem[37][3] ), .B(\u_div/PartRem[37][2] ), .Y(
        \u_div/SumTmp[36][3] ) );
  XNOR2X1 U355 ( .A(\u_div/PartRem[36][3] ), .B(\u_div/PartRem[36][2] ), .Y(
        \u_div/SumTmp[35][3] ) );
  OR2X1 U356 ( .A(\u_div/PartRem[35][5] ), .B(\u_div/u_add_PartRem_2_34/n2 ), 
        .Y(\u_div/CryTmp[34][6] ) );
  XNOR2X1 U357 ( .A(\u_div/PartRem[35][3] ), .B(\u_div/PartRem[35][2] ), .Y(
        \u_div/SumTmp[34][3] ) );
  OR2X1 U358 ( .A(\u_div/PartRem[34][5] ), .B(\u_div/u_add_PartRem_2_33/n2 ), 
        .Y(\u_div/CryTmp[33][6] ) );
  XNOR2X1 U359 ( .A(\u_div/PartRem[34][3] ), .B(\u_div/PartRem[34][2] ), .Y(
        \u_div/SumTmp[33][3] ) );
  OR2X1 U360 ( .A(\u_div/PartRem[33][5] ), .B(\u_div/u_add_PartRem_2_32/n2 ), 
        .Y(\u_div/CryTmp[32][6] ) );
  XNOR2X1 U361 ( .A(\u_div/PartRem[33][3] ), .B(\u_div/PartRem[33][2] ), .Y(
        \u_div/SumTmp[32][3] ) );
  OR2X1 U362 ( .A(\u_div/PartRem[33][2] ), .B(\u_div/PartRem[33][3] ), .Y(
        \u_div/u_add_PartRem_2_32/n3 ) );
  OR2X1 U363 ( .A(\u_div/PartRem[32][5] ), .B(\u_div/u_add_PartRem_2_31/n2 ), 
        .Y(\u_div/CryTmp[31][6] ) );
  XNOR2X1 U364 ( .A(\u_div/PartRem[32][3] ), .B(\u_div/PartRem[32][2] ), .Y(
        \u_div/SumTmp[31][3] ) );
  XNOR2X1 U365 ( .A(\u_div/PartRem[31][3] ), .B(\u_div/PartRem[31][2] ), .Y(
        \u_div/SumTmp[30][3] ) );
  XNOR2X1 U366 ( .A(\u_div/PartRem[30][3] ), .B(\u_div/PartRem[30][2] ), .Y(
        \u_div/SumTmp[29][3] ) );
  XNOR2X1 U367 ( .A(\u_div/PartRem[29][3] ), .B(\u_div/PartRem[29][2] ), .Y(
        \u_div/SumTmp[28][3] ) );
  OR2X1 U368 ( .A(\u_div/PartRem[28][5] ), .B(\u_div/u_add_PartRem_2_27/n2 ), 
        .Y(\u_div/CryTmp[27][6] ) );
  XNOR2X1 U369 ( .A(\u_div/PartRem[28][3] ), .B(\u_div/PartRem[28][2] ), .Y(
        \u_div/SumTmp[27][3] ) );
  OR2X1 U370 ( .A(\u_div/PartRem[28][2] ), .B(\u_div/PartRem[28][3] ), .Y(
        \u_div/u_add_PartRem_2_27/n3 ) );
  OR2X1 U371 ( .A(\u_div/PartRem[27][5] ), .B(\u_div/u_add_PartRem_2_26/n2 ), 
        .Y(\u_div/CryTmp[26][6] ) );
  XNOR2X1 U372 ( .A(\u_div/PartRem[27][3] ), .B(\u_div/PartRem[27][2] ), .Y(
        \u_div/SumTmp[26][3] ) );
  XNOR2X1 U373 ( .A(\u_div/PartRem[26][3] ), .B(\u_div/PartRem[26][2] ), .Y(
        \u_div/SumTmp[25][3] ) );
  OR2X1 U374 ( .A(\u_div/PartRem[25][5] ), .B(\u_div/u_add_PartRem_2_24/n2 ), 
        .Y(\u_div/CryTmp[24][6] ) );
  XNOR2X1 U375 ( .A(\u_div/PartRem[25][3] ), .B(\u_div/PartRem[25][2] ), .Y(
        \u_div/SumTmp[24][3] ) );
  OR2X1 U376 ( .A(\u_div/PartRem[24][5] ), .B(\u_div/u_add_PartRem_2_23/n2 ), 
        .Y(\u_div/CryTmp[23][6] ) );
  XNOR2X1 U377 ( .A(\u_div/PartRem[24][3] ), .B(\u_div/PartRem[24][2] ), .Y(
        \u_div/SumTmp[23][3] ) );
  OR2X1 U378 ( .A(\u_div/PartRem[23][5] ), .B(\u_div/u_add_PartRem_2_22/n2 ), 
        .Y(\u_div/CryTmp[22][6] ) );
  XNOR2X1 U379 ( .A(\u_div/PartRem[23][3] ), .B(\u_div/PartRem[23][2] ), .Y(
        \u_div/SumTmp[22][3] ) );
  OR2X1 U380 ( .A(\u_div/PartRem[23][2] ), .B(\u_div/PartRem[23][3] ), .Y(
        \u_div/u_add_PartRem_2_22/n3 ) );
  OR2X1 U381 ( .A(\u_div/PartRem[22][5] ), .B(\u_div/u_add_PartRem_2_21/n2 ), 
        .Y(\u_div/CryTmp[21][6] ) );
  XNOR2X1 U382 ( .A(\u_div/PartRem[22][3] ), .B(\u_div/PartRem[22][2] ), .Y(
        \u_div/SumTmp[21][3] ) );
  XNOR2X1 U383 ( .A(\u_div/PartRem[21][3] ), .B(\u_div/PartRem[21][2] ), .Y(
        \u_div/SumTmp[20][3] ) );
  XNOR2X1 U384 ( .A(\u_div/PartRem[20][3] ), .B(\u_div/PartRem[20][2] ), .Y(
        \u_div/SumTmp[19][3] ) );
  XNOR2X1 U385 ( .A(\u_div/PartRem[19][3] ), .B(\u_div/PartRem[19][2] ), .Y(
        \u_div/SumTmp[18][3] ) );
  OR2X1 U386 ( .A(\u_div/PartRem[18][5] ), .B(\u_div/u_add_PartRem_2_17/n2 ), 
        .Y(\u_div/CryTmp[17][6] ) );
  XNOR2X1 U387 ( .A(\u_div/PartRem[18][3] ), .B(\u_div/PartRem[18][2] ), .Y(
        \u_div/SumTmp[17][3] ) );
  OR2X1 U388 ( .A(\u_div/PartRem[18][2] ), .B(\u_div/PartRem[18][3] ), .Y(
        \u_div/u_add_PartRem_2_17/n3 ) );
  OR2X1 U389 ( .A(\u_div/PartRem[17][5] ), .B(\u_div/u_add_PartRem_2_16/n2 ), 
        .Y(\u_div/CryTmp[16][6] ) );
  XNOR2X1 U390 ( .A(\u_div/PartRem[17][3] ), .B(\u_div/PartRem[17][2] ), .Y(
        \u_div/SumTmp[16][3] ) );
  XNOR2X1 U391 ( .A(\u_div/PartRem[16][3] ), .B(\u_div/PartRem[16][2] ), .Y(
        \u_div/SumTmp[15][3] ) );
  OR2X1 U392 ( .A(\u_div/PartRem[15][5] ), .B(\u_div/u_add_PartRem_2_14/n2 ), 
        .Y(\u_div/CryTmp[14][6] ) );
  XNOR2X1 U393 ( .A(\u_div/PartRem[15][3] ), .B(\u_div/PartRem[15][2] ), .Y(
        \u_div/SumTmp[14][3] ) );
  OR2X1 U394 ( .A(\u_div/PartRem[14][5] ), .B(\u_div/u_add_PartRem_2_13/n2 ), 
        .Y(\u_div/CryTmp[13][6] ) );
  XNOR2X1 U395 ( .A(\u_div/PartRem[14][3] ), .B(\u_div/PartRem[14][2] ), .Y(
        \u_div/SumTmp[13][3] ) );
  OR2X1 U396 ( .A(\u_div/PartRem[13][5] ), .B(\u_div/u_add_PartRem_2_12/n2 ), 
        .Y(\u_div/CryTmp[12][6] ) );
  XNOR2X1 U397 ( .A(\u_div/PartRem[13][3] ), .B(\u_div/PartRem[13][2] ), .Y(
        \u_div/SumTmp[12][3] ) );
  OR2X1 U398 ( .A(\u_div/PartRem[13][2] ), .B(\u_div/PartRem[13][3] ), .Y(
        \u_div/u_add_PartRem_2_12/n3 ) );
  OR2X1 U399 ( .A(\u_div/PartRem[12][5] ), .B(\u_div/u_add_PartRem_2_11/n2 ), 
        .Y(\u_div/CryTmp[11][6] ) );
  XNOR2X1 U400 ( .A(\u_div/PartRem[12][3] ), .B(\u_div/PartRem[12][2] ), .Y(
        \u_div/SumTmp[11][3] ) );
  XNOR2X1 U401 ( .A(\u_div/PartRem[11][3] ), .B(\u_div/PartRem[11][2] ), .Y(
        \u_div/SumTmp[10][3] ) );
  XNOR2X1 U402 ( .A(\u_div/PartRem[10][3] ), .B(\u_div/PartRem[10][2] ), .Y(
        \u_div/SumTmp[9][3] ) );
  XNOR2X1 U403 ( .A(\u_div/PartRem[9][3] ), .B(\u_div/PartRem[9][2] ), .Y(
        \u_div/SumTmp[8][3] ) );
  XNOR2X1 U404 ( .A(\u_div/PartRem[8][3] ), .B(\u_div/PartRem[8][2] ), .Y(
        \u_div/SumTmp[7][3] ) );
  OR2X1 U405 ( .A(\u_div/PartRem[8][2] ), .B(\u_div/PartRem[8][3] ), .Y(
        \u_div/u_add_PartRem_2_7/n3 ) );
  XNOR2X1 U406 ( .A(\u_div/PartRem[7][3] ), .B(\u_div/PartRem[7][2] ), .Y(
        \u_div/SumTmp[6][3] ) );
  XNOR2X1 U407 ( .A(\u_div/PartRem[6][3] ), .B(\u_div/PartRem[6][2] ), .Y(
        \u_div/SumTmp[5][3] ) );
  XNOR2X1 U408 ( .A(\u_div/PartRem[5][3] ), .B(\u_div/PartRem[5][2] ), .Y(
        \u_div/SumTmp[4][3] ) );
  XNOR2X1 U409 ( .A(\u_div/PartRem[4][3] ), .B(\u_div/PartRem[4][2] ), .Y(
        \u_div/SumTmp[3][3] ) );
  XNOR2X1 U410 ( .A(\u_div/PartRem[3][3] ), .B(\u_div/PartRem[3][2] ), .Y(
        \u_div/SumTmp[2][3] ) );
  OR2X1 U411 ( .A(\u_div/PartRem[3][2] ), .B(\u_div/PartRem[3][3] ), .Y(
        \u_div/u_add_PartRem_2_2/n3 ) );
  OR2X1 U412 ( .A(\u_div/PartRem[2][5] ), .B(\u_div/u_add_PartRem_2_1/n2 ), 
        .Y(\u_div/CryTmp[1][6] ) );
  XNOR2X1 U413 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/PartRem[2][2] ), .Y(
        \u_div/SumTmp[1][3] ) );
  NAND2BX1 U414 ( .AN(\u_div/PartRem[1][3] ), .B(n1), .Y(n6) );
  XNOR2X1 U415 ( .A(\u_div/PartRem[63][0] ), .B(\u_div/PartRem[62][0] ), .Y(
        \u_div/SumTmp[59][3] ) );
  XOR2X1 U416 ( .A(\u_div/CryTmp[58][6] ), .B(n4), .Y(\u_div/QInv[58] ) );
  XOR2X1 U417 ( .A(\u_div/CryTmp[39][6] ), .B(n4), .Y(\u_div/QInv[39] ) );
  XOR2X1 U418 ( .A(\u_div/CryTmp[29][6] ), .B(n4), .Y(\u_div/QInv[29] ) );
  XOR2X1 U419 ( .A(\u_div/CryTmp[18][6] ), .B(n4), .Y(\u_div/QInv[18] ) );
  XOR2X1 U420 ( .A(\u_div/CryTmp[0][6] ), .B(n4), .Y(\u_div/QInv[0] ) );
endmodule


module GSIM_DW01_inc_3 ( A, SUM );
  input [63:0] A;
  output [63:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;

  NOR3BX1 U2 ( .AN(A[59]), .B(n1), .C(n24), .Y(n22) );
  XOR2X1 U3 ( .A(A[63]), .B(n20), .Y(SUM[63]) );
  NOR2BX1 U4 ( .AN(A[62]), .B(n21), .Y(n20) );
  NOR3BX1 U5 ( .AN(A[55]), .B(n2), .C(n30), .Y(n28) );
  XNOR2X1 U6 ( .A(A[62]), .B(n21), .Y(SUM[62]) );
  NOR3BX1 U7 ( .AN(A[51]), .B(n3), .C(n34), .Y(n32) );
  NOR3BX1 U8 ( .AN(A[47]), .B(n4), .C(n38), .Y(n36) );
  NOR3BX1 U9 ( .AN(A[43]), .B(n5), .C(n42), .Y(n40) );
  NOR3BX1 U10 ( .AN(A[39]), .B(n6), .C(n46), .Y(n44) );
  NOR3BX1 U11 ( .AN(A[35]), .B(n7), .C(n52), .Y(n50) );
  NOR3BX1 U12 ( .AN(A[31]), .B(n8), .C(n56), .Y(n54) );
  NOR3BX1 U13 ( .AN(A[27]), .B(n9), .C(n60), .Y(n58) );
  NOR3BX1 U14 ( .AN(A[23]), .B(n10), .C(n64), .Y(n62) );
  NOR3BX1 U15 ( .AN(A[19]), .B(n11), .C(n68), .Y(n66) );
  NOR3BX1 U16 ( .AN(A[15]), .B(n12), .C(n72), .Y(n70) );
  NOR3BX1 U17 ( .AN(A[11]), .B(n13), .C(n76), .Y(n74) );
  NOR3BX1 U18 ( .AN(A[7]), .B(n14), .C(n19), .Y(n17) );
  NAND3X1 U19 ( .A(A[4]), .B(n26), .C(A[5]), .Y(n19) );
  NOR3BX1 U20 ( .AN(A[3]), .B(n15), .C(n48), .Y(n26) );
  NOR2XL U21 ( .A(n24), .B(n1), .Y(n27) );
  NAND2XL U22 ( .A(A[56]), .B(n28), .Y(n29) );
  NOR2XL U23 ( .A(n30), .B(n2), .Y(n31) );
  NAND2XL U24 ( .A(A[52]), .B(n32), .Y(n33) );
  NOR2XL U25 ( .A(n34), .B(n3), .Y(n35) );
  NAND2XL U26 ( .A(A[48]), .B(n36), .Y(n37) );
  NOR2XL U27 ( .A(n38), .B(n4), .Y(n39) );
  NAND2XL U28 ( .A(A[44]), .B(n40), .Y(n41) );
  NOR2XL U29 ( .A(n42), .B(n5), .Y(n43) );
  NAND2XL U30 ( .A(A[40]), .B(n44), .Y(n45) );
  NOR2XL U31 ( .A(n46), .B(n6), .Y(n49) );
  NAND2XL U32 ( .A(A[36]), .B(n50), .Y(n51) );
  NOR2XL U33 ( .A(n52), .B(n7), .Y(n53) );
  NAND2XL U34 ( .A(A[32]), .B(n54), .Y(n55) );
  NOR2XL U35 ( .A(n56), .B(n8), .Y(n57) );
  NAND2XL U36 ( .A(A[28]), .B(n58), .Y(n59) );
  NOR2XL U37 ( .A(n60), .B(n9), .Y(n61) );
  NAND2XL U38 ( .A(A[24]), .B(n62), .Y(n63) );
  NOR2XL U39 ( .A(n64), .B(n10), .Y(n65) );
  NAND2XL U40 ( .A(A[20]), .B(n66), .Y(n67) );
  NOR2XL U41 ( .A(n68), .B(n11), .Y(n69) );
  NAND2XL U42 ( .A(A[16]), .B(n70), .Y(n71) );
  NOR2XL U43 ( .A(n72), .B(n12), .Y(n73) );
  NAND2XL U44 ( .A(A[12]), .B(n74), .Y(n75) );
  NOR2XL U45 ( .A(n76), .B(n13), .Y(n77) );
  NAND2XL U46 ( .A(A[8]), .B(n17), .Y(n16) );
  NOR2XL U47 ( .A(n19), .B(n14), .Y(n18) );
  NAND2XL U48 ( .A(A[4]), .B(n26), .Y(n25) );
  XOR2XL U49 ( .A(A[60]), .B(n22), .Y(SUM[60]) );
  NAND2XL U50 ( .A(A[60]), .B(n22), .Y(n23) );
  NOR2XL U51 ( .A(n48), .B(n15), .Y(n47) );
  CLKINVX1 U52 ( .A(A[58]), .Y(n1) );
  CLKINVX1 U53 ( .A(A[54]), .Y(n2) );
  CLKINVX1 U54 ( .A(A[50]), .Y(n3) );
  CLKINVX1 U55 ( .A(A[46]), .Y(n4) );
  CLKINVX1 U56 ( .A(A[42]), .Y(n5) );
  CLKINVX1 U57 ( .A(A[38]), .Y(n6) );
  CLKINVX1 U58 ( .A(A[34]), .Y(n7) );
  CLKINVX1 U59 ( .A(A[30]), .Y(n8) );
  CLKINVX1 U60 ( .A(A[2]), .Y(n15) );
  CLKINVX1 U61 ( .A(A[26]), .Y(n9) );
  CLKINVX1 U62 ( .A(A[22]), .Y(n10) );
  CLKINVX1 U63 ( .A(A[14]), .Y(n12) );
  CLKINVX1 U64 ( .A(A[10]), .Y(n13) );
  CLKINVX1 U65 ( .A(A[6]), .Y(n14) );
  CLKINVX1 U66 ( .A(A[18]), .Y(n11) );
  XNOR2X1 U67 ( .A(A[9]), .B(n16), .Y(SUM[9]) );
  XOR2X1 U68 ( .A(A[8]), .B(n17), .Y(SUM[8]) );
  XOR2X1 U69 ( .A(A[7]), .B(n18), .Y(SUM[7]) );
  XOR2X1 U70 ( .A(n14), .B(n19), .Y(SUM[6]) );
  NAND3X1 U71 ( .A(A[60]), .B(n22), .C(A[61]), .Y(n21) );
  XNOR2X1 U72 ( .A(A[61]), .B(n23), .Y(SUM[61]) );
  XNOR2X1 U73 ( .A(A[5]), .B(n25), .Y(SUM[5]) );
  XOR2X1 U74 ( .A(A[59]), .B(n27), .Y(SUM[59]) );
  XOR2X1 U75 ( .A(n1), .B(n24), .Y(SUM[58]) );
  NAND3X1 U76 ( .A(A[56]), .B(n28), .C(A[57]), .Y(n24) );
  XNOR2X1 U77 ( .A(A[57]), .B(n29), .Y(SUM[57]) );
  XOR2X1 U78 ( .A(A[56]), .B(n28), .Y(SUM[56]) );
  XOR2X1 U79 ( .A(A[55]), .B(n31), .Y(SUM[55]) );
  XOR2X1 U80 ( .A(n2), .B(n30), .Y(SUM[54]) );
  NAND3X1 U81 ( .A(A[52]), .B(n32), .C(A[53]), .Y(n30) );
  XNOR2X1 U82 ( .A(A[53]), .B(n33), .Y(SUM[53]) );
  XOR2X1 U83 ( .A(A[52]), .B(n32), .Y(SUM[52]) );
  XOR2X1 U84 ( .A(A[51]), .B(n35), .Y(SUM[51]) );
  XOR2X1 U85 ( .A(n3), .B(n34), .Y(SUM[50]) );
  NAND3X1 U86 ( .A(A[48]), .B(n36), .C(A[49]), .Y(n34) );
  XOR2X1 U87 ( .A(A[4]), .B(n26), .Y(SUM[4]) );
  XNOR2X1 U88 ( .A(A[49]), .B(n37), .Y(SUM[49]) );
  XOR2X1 U89 ( .A(A[48]), .B(n36), .Y(SUM[48]) );
  XOR2X1 U90 ( .A(A[47]), .B(n39), .Y(SUM[47]) );
  XOR2X1 U91 ( .A(n4), .B(n38), .Y(SUM[46]) );
  NAND3X1 U92 ( .A(A[44]), .B(n40), .C(A[45]), .Y(n38) );
  XNOR2X1 U93 ( .A(A[45]), .B(n41), .Y(SUM[45]) );
  XOR2X1 U94 ( .A(A[44]), .B(n40), .Y(SUM[44]) );
  XOR2X1 U95 ( .A(A[43]), .B(n43), .Y(SUM[43]) );
  XOR2X1 U96 ( .A(n5), .B(n42), .Y(SUM[42]) );
  NAND3X1 U97 ( .A(A[40]), .B(n44), .C(A[41]), .Y(n42) );
  XNOR2X1 U98 ( .A(A[41]), .B(n45), .Y(SUM[41]) );
  XOR2X1 U99 ( .A(A[40]), .B(n44), .Y(SUM[40]) );
  XOR2X1 U100 ( .A(A[3]), .B(n47), .Y(SUM[3]) );
  XOR2X1 U101 ( .A(A[39]), .B(n49), .Y(SUM[39]) );
  XOR2X1 U102 ( .A(n6), .B(n46), .Y(SUM[38]) );
  NAND3X1 U103 ( .A(A[36]), .B(n50), .C(A[37]), .Y(n46) );
  XNOR2X1 U104 ( .A(A[37]), .B(n51), .Y(SUM[37]) );
  XOR2X1 U105 ( .A(A[36]), .B(n50), .Y(SUM[36]) );
  XOR2X1 U106 ( .A(A[35]), .B(n53), .Y(SUM[35]) );
  XOR2X1 U107 ( .A(n7), .B(n52), .Y(SUM[34]) );
  NAND3X1 U108 ( .A(A[32]), .B(n54), .C(A[33]), .Y(n52) );
  XNOR2X1 U109 ( .A(A[33]), .B(n55), .Y(SUM[33]) );
  XOR2X1 U110 ( .A(A[32]), .B(n54), .Y(SUM[32]) );
  XOR2X1 U111 ( .A(A[31]), .B(n57), .Y(SUM[31]) );
  XOR2X1 U112 ( .A(n8), .B(n56), .Y(SUM[30]) );
  NAND3X1 U113 ( .A(A[28]), .B(n58), .C(A[29]), .Y(n56) );
  XOR2X1 U114 ( .A(n15), .B(n48), .Y(SUM[2]) );
  XNOR2X1 U115 ( .A(A[29]), .B(n59), .Y(SUM[29]) );
  XOR2X1 U116 ( .A(A[28]), .B(n58), .Y(SUM[28]) );
  XOR2X1 U117 ( .A(A[27]), .B(n61), .Y(SUM[27]) );
  XOR2X1 U118 ( .A(n9), .B(n60), .Y(SUM[26]) );
  NAND3X1 U119 ( .A(A[24]), .B(n62), .C(A[25]), .Y(n60) );
  XNOR2X1 U120 ( .A(A[25]), .B(n63), .Y(SUM[25]) );
  XOR2X1 U121 ( .A(A[24]), .B(n62), .Y(SUM[24]) );
  XOR2X1 U122 ( .A(A[23]), .B(n65), .Y(SUM[23]) );
  XOR2X1 U123 ( .A(n10), .B(n64), .Y(SUM[22]) );
  NAND3X1 U124 ( .A(A[20]), .B(n66), .C(A[21]), .Y(n64) );
  XNOR2X1 U125 ( .A(A[21]), .B(n67), .Y(SUM[21]) );
  XOR2X1 U126 ( .A(A[20]), .B(n66), .Y(SUM[20]) );
  XOR2X1 U127 ( .A(A[19]), .B(n69), .Y(SUM[19]) );
  XOR2X1 U128 ( .A(n11), .B(n68), .Y(SUM[18]) );
  NAND3X1 U129 ( .A(A[16]), .B(n70), .C(A[17]), .Y(n68) );
  XNOR2X1 U130 ( .A(A[17]), .B(n71), .Y(SUM[17]) );
  XOR2X1 U131 ( .A(A[16]), .B(n70), .Y(SUM[16]) );
  XOR2X1 U132 ( .A(A[15]), .B(n73), .Y(SUM[15]) );
  XOR2X1 U133 ( .A(n12), .B(n72), .Y(SUM[14]) );
  NAND3X1 U134 ( .A(A[12]), .B(n74), .C(A[13]), .Y(n72) );
  XNOR2X1 U135 ( .A(A[13]), .B(n75), .Y(SUM[13]) );
  XOR2X1 U136 ( .A(A[12]), .B(n74), .Y(SUM[12]) );
  XOR2X1 U137 ( .A(A[11]), .B(n77), .Y(SUM[11]) );
  XOR2X1 U138 ( .A(n13), .B(n76), .Y(SUM[10]) );
  NAND3X1 U139 ( .A(A[8]), .B(n17), .C(A[9]), .Y(n76) );
  NAND2X1 U140 ( .A(A[1]), .B(A[0]), .Y(n48) );
endmodule


module GSIM_DW01_absval_1 ( A, ABSVAL );
  input [63:0] A;
  output [63:0] ABSVAL;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68;
  wire   [63:0] AMUX1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  GSIM_DW01_inc_3 NEG ( .A({n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
        n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
        n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
        n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
        n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68}), .SUM({
        AMUX1[63:2], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1}) );
  CLKINVX1 U1 ( .A(A[61]), .Y(n7) );
  CLKMX2X2 U2 ( .A(A[61]), .B(AMUX1[61]), .S0(n4), .Y(ABSVAL[61]) );
  CLKINVX1 U3 ( .A(A[3]), .Y(n65) );
  INVX3 U4 ( .A(n5), .Y(n4) );
  INVX3 U5 ( .A(n5), .Y(n3) );
  INVX3 U6 ( .A(n5), .Y(n2) );
  INVX3 U7 ( .A(n5), .Y(n1) );
  CLKINVX1 U8 ( .A(A[63]), .Y(n5) );
  CLKINVX1 U9 ( .A(A[58]), .Y(n10) );
  CLKINVX1 U10 ( .A(A[62]), .Y(n6) );
  CLKINVX1 U11 ( .A(A[59]), .Y(n9) );
  CLKINVX1 U12 ( .A(A[55]), .Y(n13) );
  CLKINVX1 U13 ( .A(A[51]), .Y(n17) );
  CLKINVX1 U14 ( .A(A[47]), .Y(n21) );
  CLKINVX1 U15 ( .A(A[60]), .Y(n8) );
  CLKINVX1 U16 ( .A(A[56]), .Y(n12) );
  CLKINVX1 U17 ( .A(A[52]), .Y(n16) );
  CLKINVX1 U18 ( .A(A[48]), .Y(n20) );
  CLKINVX1 U19 ( .A(A[54]), .Y(n14) );
  CLKINVX1 U20 ( .A(A[50]), .Y(n18) );
  CLKINVX1 U21 ( .A(A[46]), .Y(n22) );
  CLKINVX1 U22 ( .A(A[42]), .Y(n26) );
  CLKINVX1 U23 ( .A(A[38]), .Y(n30) );
  CLKINVX1 U24 ( .A(A[34]), .Y(n34) );
  CLKINVX1 U25 ( .A(A[30]), .Y(n38) );
  CLKINVX1 U26 ( .A(A[2]), .Y(n66) );
  CLKINVX1 U27 ( .A(A[57]), .Y(n11) );
  CLKINVX1 U28 ( .A(A[53]), .Y(n15) );
  CLKINVX1 U29 ( .A(A[49]), .Y(n19) );
  CLKINVX1 U30 ( .A(A[45]), .Y(n23) );
  CLKINVX1 U31 ( .A(A[41]), .Y(n27) );
  CLKINVX1 U32 ( .A(A[37]), .Y(n31) );
  CLKINVX1 U33 ( .A(A[33]), .Y(n35) );
  CLKINVX1 U34 ( .A(A[43]), .Y(n25) );
  CLKINVX1 U35 ( .A(A[39]), .Y(n29) );
  CLKINVX1 U36 ( .A(A[35]), .Y(n33) );
  CLKINVX1 U37 ( .A(A[31]), .Y(n37) );
  CLKINVX1 U38 ( .A(A[27]), .Y(n41) );
  CLKINVX1 U39 ( .A(A[23]), .Y(n45) );
  CLKINVX1 U40 ( .A(A[19]), .Y(n49) );
  CLKINVX1 U41 ( .A(A[15]), .Y(n53) );
  CLKINVX1 U42 ( .A(A[44]), .Y(n24) );
  CLKINVX1 U43 ( .A(A[40]), .Y(n28) );
  CLKINVX1 U44 ( .A(A[36]), .Y(n32) );
  CLKINVX1 U45 ( .A(A[32]), .Y(n36) );
  CLKINVX1 U46 ( .A(A[28]), .Y(n40) );
  CLKINVX1 U47 ( .A(A[24]), .Y(n44) );
  CLKINVX1 U48 ( .A(A[20]), .Y(n48) );
  CLKINVX1 U49 ( .A(A[16]), .Y(n52) );
  CLKINVX1 U50 ( .A(A[4]), .Y(n64) );
  CLKINVX1 U51 ( .A(A[26]), .Y(n42) );
  CLKINVX1 U52 ( .A(A[22]), .Y(n46) );
  CLKINVX1 U53 ( .A(A[14]), .Y(n54) );
  CLKINVX1 U54 ( .A(A[10]), .Y(n58) );
  CLKINVX1 U55 ( .A(A[6]), .Y(n62) );
  CLKINVX1 U56 ( .A(A[29]), .Y(n39) );
  CLKINVX1 U57 ( .A(A[25]), .Y(n43) );
  CLKINVX1 U58 ( .A(A[21]), .Y(n47) );
  CLKINVX1 U59 ( .A(A[17]), .Y(n51) );
  CLKINVX1 U60 ( .A(A[13]), .Y(n55) );
  CLKINVX1 U61 ( .A(A[9]), .Y(n59) );
  CLKINVX1 U62 ( .A(A[5]), .Y(n63) );
  CLKINVX1 U63 ( .A(A[11]), .Y(n57) );
  CLKINVX1 U64 ( .A(A[7]), .Y(n61) );
  CLKINVX1 U65 ( .A(A[18]), .Y(n50) );
  CLKINVX1 U66 ( .A(A[12]), .Y(n56) );
  CLKINVX1 U67 ( .A(A[8]), .Y(n60) );
  CLKINVX1 U68 ( .A(A[0]), .Y(n68) );
  CLKINVX1 U69 ( .A(A[1]), .Y(n67) );
  CLKMX2X2 U70 ( .A(A[9]), .B(AMUX1[9]), .S0(n3), .Y(ABSVAL[9]) );
  CLKMX2X2 U71 ( .A(A[8]), .B(AMUX1[8]), .S0(n4), .Y(ABSVAL[8]) );
  CLKMX2X2 U72 ( .A(A[7]), .B(AMUX1[7]), .S0(n4), .Y(ABSVAL[7]) );
  CLKMX2X2 U73 ( .A(A[6]), .B(AMUX1[6]), .S0(n4), .Y(ABSVAL[6]) );
  AND2X1 U74 ( .A(AMUX1[63]), .B(n4), .Y(ABSVAL[63]) );
  CLKMX2X2 U75 ( .A(A[62]), .B(AMUX1[62]), .S0(n4), .Y(ABSVAL[62]) );
  CLKMX2X2 U76 ( .A(A[60]), .B(AMUX1[60]), .S0(n4), .Y(ABSVAL[60]) );
  CLKMX2X2 U77 ( .A(A[5]), .B(AMUX1[5]), .S0(n4), .Y(ABSVAL[5]) );
  CLKMX2X2 U78 ( .A(A[59]), .B(AMUX1[59]), .S0(n4), .Y(ABSVAL[59]) );
  CLKMX2X2 U79 ( .A(A[58]), .B(AMUX1[58]), .S0(n4), .Y(ABSVAL[58]) );
  CLKMX2X2 U80 ( .A(A[57]), .B(AMUX1[57]), .S0(n4), .Y(ABSVAL[57]) );
  CLKMX2X2 U81 ( .A(A[56]), .B(AMUX1[56]), .S0(n3), .Y(ABSVAL[56]) );
  CLKMX2X2 U82 ( .A(A[55]), .B(AMUX1[55]), .S0(n3), .Y(ABSVAL[55]) );
  CLKMX2X2 U83 ( .A(A[54]), .B(AMUX1[54]), .S0(n3), .Y(ABSVAL[54]) );
  CLKMX2X2 U84 ( .A(A[53]), .B(AMUX1[53]), .S0(n3), .Y(ABSVAL[53]) );
  CLKMX2X2 U85 ( .A(A[52]), .B(AMUX1[52]), .S0(n3), .Y(ABSVAL[52]) );
  CLKMX2X2 U86 ( .A(A[51]), .B(AMUX1[51]), .S0(n3), .Y(ABSVAL[51]) );
  CLKMX2X2 U87 ( .A(A[50]), .B(AMUX1[50]), .S0(n3), .Y(ABSVAL[50]) );
  CLKMX2X2 U88 ( .A(A[4]), .B(AMUX1[4]), .S0(n3), .Y(ABSVAL[4]) );
  CLKMX2X2 U89 ( .A(A[49]), .B(AMUX1[49]), .S0(n3), .Y(ABSVAL[49]) );
  CLKMX2X2 U90 ( .A(A[48]), .B(AMUX1[48]), .S0(n3), .Y(ABSVAL[48]) );
  CLKMX2X2 U91 ( .A(A[47]), .B(AMUX1[47]), .S0(n3), .Y(ABSVAL[47]) );
  CLKMX2X2 U92 ( .A(A[46]), .B(AMUX1[46]), .S0(n3), .Y(ABSVAL[46]) );
  CLKMX2X2 U93 ( .A(A[45]), .B(AMUX1[45]), .S0(n3), .Y(ABSVAL[45]) );
  CLKMX2X2 U94 ( .A(A[44]), .B(AMUX1[44]), .S0(n2), .Y(ABSVAL[44]) );
  CLKMX2X2 U95 ( .A(A[43]), .B(AMUX1[43]), .S0(n2), .Y(ABSVAL[43]) );
  CLKMX2X2 U96 ( .A(A[42]), .B(AMUX1[42]), .S0(n2), .Y(ABSVAL[42]) );
  CLKMX2X2 U97 ( .A(A[41]), .B(AMUX1[41]), .S0(n2), .Y(ABSVAL[41]) );
  CLKMX2X2 U98 ( .A(A[40]), .B(AMUX1[40]), .S0(n2), .Y(ABSVAL[40]) );
  CLKMX2X2 U99 ( .A(A[3]), .B(AMUX1[3]), .S0(n2), .Y(ABSVAL[3]) );
  CLKMX2X2 U100 ( .A(A[39]), .B(AMUX1[39]), .S0(n2), .Y(ABSVAL[39]) );
  CLKMX2X2 U101 ( .A(A[38]), .B(AMUX1[38]), .S0(n2), .Y(ABSVAL[38]) );
  CLKMX2X2 U102 ( .A(A[37]), .B(AMUX1[37]), .S0(n2), .Y(ABSVAL[37]) );
  CLKMX2X2 U103 ( .A(A[36]), .B(AMUX1[36]), .S0(n2), .Y(ABSVAL[36]) );
  CLKMX2X2 U104 ( .A(A[35]), .B(AMUX1[35]), .S0(n2), .Y(ABSVAL[35]) );
  CLKMX2X2 U105 ( .A(A[34]), .B(AMUX1[34]), .S0(n2), .Y(ABSVAL[34]) );
  CLKMX2X2 U106 ( .A(A[33]), .B(AMUX1[33]), .S0(n1), .Y(ABSVAL[33]) );
  CLKMX2X2 U107 ( .A(A[32]), .B(AMUX1[32]), .S0(n1), .Y(ABSVAL[32]) );
  CLKMX2X2 U108 ( .A(A[31]), .B(AMUX1[31]), .S0(n1), .Y(ABSVAL[31]) );
  CLKMX2X2 U109 ( .A(A[30]), .B(AMUX1[30]), .S0(n1), .Y(ABSVAL[30]) );
  CLKMX2X2 U110 ( .A(A[2]), .B(AMUX1[2]), .S0(n1), .Y(ABSVAL[2]) );
  CLKMX2X2 U111 ( .A(A[29]), .B(AMUX1[29]), .S0(n1), .Y(ABSVAL[29]) );
  CLKMX2X2 U112 ( .A(A[28]), .B(AMUX1[28]), .S0(n1), .Y(ABSVAL[28]) );
  CLKMX2X2 U113 ( .A(A[27]), .B(AMUX1[27]), .S0(n1), .Y(ABSVAL[27]) );
  CLKMX2X2 U114 ( .A(A[26]), .B(AMUX1[26]), .S0(n1), .Y(ABSVAL[26]) );
  CLKMX2X2 U115 ( .A(A[25]), .B(AMUX1[25]), .S0(n1), .Y(ABSVAL[25]) );
  CLKMX2X2 U116 ( .A(A[24]), .B(AMUX1[24]), .S0(n1), .Y(ABSVAL[24]) );
  CLKMX2X2 U117 ( .A(A[23]), .B(AMUX1[23]), .S0(n1), .Y(ABSVAL[23]) );
  CLKMX2X2 U118 ( .A(A[22]), .B(AMUX1[22]), .S0(n1), .Y(ABSVAL[22]) );
  CLKMX2X2 U119 ( .A(A[21]), .B(AMUX1[21]), .S0(n1), .Y(ABSVAL[21]) );
  CLKMX2X2 U120 ( .A(A[20]), .B(AMUX1[20]), .S0(n1), .Y(ABSVAL[20]) );
  CLKMX2X2 U121 ( .A(A[19]), .B(AMUX1[19]), .S0(n1), .Y(ABSVAL[19]) );
  CLKMX2X2 U122 ( .A(A[18]), .B(AMUX1[18]), .S0(n1), .Y(ABSVAL[18]) );
  CLKMX2X2 U123 ( .A(A[17]), .B(AMUX1[17]), .S0(n2), .Y(ABSVAL[17]) );
  CLKMX2X2 U124 ( .A(A[16]), .B(AMUX1[16]), .S0(n2), .Y(ABSVAL[16]) );
  CLKMX2X2 U125 ( .A(A[15]), .B(AMUX1[15]), .S0(n2), .Y(ABSVAL[15]) );
  CLKMX2X2 U126 ( .A(A[14]), .B(AMUX1[14]), .S0(n2), .Y(ABSVAL[14]) );
  CLKMX2X2 U127 ( .A(A[13]), .B(AMUX1[13]), .S0(n3), .Y(ABSVAL[13]) );
  CLKMX2X2 U128 ( .A(A[12]), .B(AMUX1[12]), .S0(n3), .Y(ABSVAL[12]) );
  CLKMX2X2 U129 ( .A(A[11]), .B(AMUX1[11]), .S0(n3), .Y(ABSVAL[11]) );
  CLKMX2X2 U130 ( .A(A[10]), .B(AMUX1[10]), .S0(n2), .Y(ABSVAL[10]) );
endmodule


module GSIM_DW_inc_1 ( carry_in, a, carry_out, sum );
  input [63:0] a;
  output [63:0] sum;
  input carry_in;
  output carry_out;
  wire   \sum[63] , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63;
  assign sum[62] = \sum[63] ;
  assign sum[61] = \sum[63] ;
  assign sum[63] = \sum[63] ;

  ADDHXL U15 ( .A(a[51]), .B(n13), .CO(n12), .S(sum[51]) );
  ADDHXL U44 ( .A(a[22]), .B(n42), .CO(n41), .S(sum[22]) );
  ADDHXL U66 ( .A(carry_in), .B(a[0]), .CO(n63), .S(sum[0]) );
  ADDHX1 U70 ( .A(a[5]), .B(n59), .CO(n58), .S(sum[5]) );
  ADDHX1 U71 ( .A(a[50]), .B(n14), .CO(n13), .S(sum[50]) );
  ADDHX1 U72 ( .A(a[58]), .B(n6), .CO(n5), .S(sum[58]) );
  XOR2X1 U73 ( .A(n4), .B(a[60]), .Y(sum[60]) );
  ADDHX2 U74 ( .A(a[3]), .B(n61), .CO(n60), .S(sum[3]) );
  ADDHX2 U75 ( .A(a[41]), .B(n23), .CO(n22), .S(sum[41]) );
  ADDHX2 U76 ( .A(a[8]), .B(n56), .CO(n55), .S(sum[8]) );
  ADDHX2 U77 ( .A(a[23]), .B(n41), .CO(n40), .S(sum[23]) );
  ADDHX2 U78 ( .A(a[18]), .B(n46), .CO(n45), .S(sum[18]) );
  ADDHX2 U79 ( .A(a[36]), .B(n28), .CO(n27), .S(sum[36]) );
  ADDHX2 U80 ( .A(a[26]), .B(n38), .CO(n37), .S(sum[26]) );
  ADDHX2 U81 ( .A(a[39]), .B(n25), .CO(n24), .S(sum[39]) );
  ADDHX2 U82 ( .A(a[34]), .B(n30), .CO(n29), .S(sum[34]) );
  ADDHX2 U83 ( .A(a[29]), .B(n35), .CO(n34), .S(sum[29]) );
  ADDHX2 U84 ( .A(a[16]), .B(n48), .CO(n47), .S(sum[16]) );
  ADDHX2 U85 ( .A(a[14]), .B(n50), .CO(n49), .S(sum[14]) );
  ADDHX2 U86 ( .A(a[31]), .B(n33), .CO(n32), .S(sum[31]) );
  ADDHX1 U87 ( .A(a[11]), .B(n53), .CO(n52), .S(sum[11]) );
  ADDHX2 U88 ( .A(a[55]), .B(n9), .CO(n8), .S(sum[55]) );
  ADDHX2 U89 ( .A(a[47]), .B(n17), .CO(n16), .S(sum[47]) );
  ADDHX2 U90 ( .A(a[44]), .B(n20), .CO(n19), .S(sum[44]) );
  ADDHXL U91 ( .A(a[12]), .B(n52), .CO(n51), .S(sum[12]) );
  ADDHXL U92 ( .A(a[4]), .B(n60), .CO(n59), .S(sum[4]) );
  ADDHX2 U93 ( .A(a[40]), .B(n24), .CO(n23), .S(sum[40]) );
  ADDHX2 U94 ( .A(a[35]), .B(n29), .CO(n28), .S(sum[35]) );
  ADDHX2 U95 ( .A(a[30]), .B(n34), .CO(n33), .S(sum[30]) );
  ADDHX2 U96 ( .A(a[13]), .B(n51), .CO(n50), .S(sum[13]) );
  ADDHX2 U97 ( .A(a[15]), .B(n49), .CO(n48), .S(sum[15]) );
  ADDHX2 U98 ( .A(a[17]), .B(n47), .CO(n46), .S(sum[17]) );
  ADDHX2 U99 ( .A(a[9]), .B(n55), .CO(n54), .S(sum[9]) );
  ADDHX2 U100 ( .A(a[37]), .B(n27), .CO(n26), .S(sum[37]) );
  ADDHX2 U101 ( .A(a[19]), .B(n45), .CO(n44), .S(sum[19]) );
  ADDHX2 U102 ( .A(a[27]), .B(n37), .CO(n36), .S(sum[27]) );
  ADDHX2 U103 ( .A(a[24]), .B(n40), .CO(n39), .S(sum[24]) );
  NOR2BX1 U104 ( .AN(a[60]), .B(n4), .Y(\sum[63] ) );
  ADDHX1 U105 ( .A(a[52]), .B(n12), .CO(n11), .S(sum[52]) );
  ADDHX1 U106 ( .A(a[1]), .B(n63), .CO(n62), .S(sum[1]) );
  ADDHX1 U107 ( .A(a[7]), .B(n57), .CO(n56), .S(sum[7]) );
  ADDHX2 U108 ( .A(a[56]), .B(n8), .CO(n7), .S(sum[56]) );
  ADDHX2 U109 ( .A(a[53]), .B(n11), .CO(n10), .S(sum[53]) );
  ADDHX2 U110 ( .A(a[48]), .B(n16), .CO(n15), .S(sum[48]) );
  ADDHX2 U111 ( .A(a[45]), .B(n19), .CO(n18), .S(sum[45]) );
  ADDHX2 U112 ( .A(a[42]), .B(n22), .CO(n21), .S(sum[42]) );
  ADDHX1 U113 ( .A(a[32]), .B(n32), .CO(n31), .S(sum[32]) );
  ADDHX1 U114 ( .A(a[21]), .B(n43), .CO(n42), .S(sum[21]) );
  ADDHX1 U115 ( .A(a[2]), .B(n62), .CO(n61), .S(sum[2]) );
  ADDHXL U116 ( .A(a[54]), .B(n10), .CO(n9), .S(sum[54]) );
  ADDHXL U117 ( .A(a[33]), .B(n31), .CO(n30), .S(sum[33]) );
  ADDHXL U118 ( .A(a[43]), .B(n21), .CO(n20), .S(sum[43]) );
  ADDHXL U119 ( .A(a[25]), .B(n39), .CO(n38), .S(sum[25]) );
  ADDHXL U120 ( .A(a[28]), .B(n36), .CO(n35), .S(sum[28]) );
  ADDHXL U121 ( .A(a[38]), .B(n26), .CO(n25), .S(sum[38]) );
  ADDHXL U122 ( .A(a[57]), .B(n7), .CO(n6), .S(sum[57]) );
  ADDHXL U123 ( .A(a[59]), .B(n5), .CO(n4), .S(sum[59]) );
  ADDHXL U124 ( .A(a[10]), .B(n54), .CO(n53), .S(sum[10]) );
  ADDHXL U125 ( .A(a[20]), .B(n44), .CO(n43), .S(sum[20]) );
  ADDHXL U126 ( .A(a[6]), .B(n58), .CO(n57), .S(sum[6]) );
  ADDHXL U127 ( .A(a[46]), .B(n18), .CO(n17), .S(sum[46]) );
  ADDHXL U128 ( .A(a[49]), .B(n15), .CO(n14), .S(sum[49]) );
endmodule


module GSIM_DW_div_tc_1 ( a, b, quotient, remainder, divide_by_0 );
  input [63:0] a;
  input [5:0] b;
  output [63:0] quotient;
  output [5:0] remainder;
  output divide_by_0;
  wire   \u_div/QInv[63] , \u_div/QInv[59] , \u_div/QInv[58] ,
         \u_div/QInv[57] , \u_div/QInv[56] , \u_div/QInv[55] ,
         \u_div/QInv[54] , \u_div/QInv[53] , \u_div/QInv[52] ,
         \u_div/QInv[51] , \u_div/QInv[50] , \u_div/QInv[49] ,
         \u_div/QInv[48] , \u_div/QInv[47] , \u_div/QInv[46] ,
         \u_div/QInv[45] , \u_div/QInv[44] , \u_div/QInv[43] ,
         \u_div/QInv[42] , \u_div/QInv[41] , \u_div/QInv[40] ,
         \u_div/QInv[39] , \u_div/QInv[38] , \u_div/QInv[37] ,
         \u_div/QInv[36] , \u_div/QInv[35] , \u_div/QInv[34] ,
         \u_div/QInv[33] , \u_div/QInv[32] , \u_div/QInv[31] ,
         \u_div/QInv[30] , \u_div/QInv[29] , \u_div/QInv[28] ,
         \u_div/QInv[27] , \u_div/QInv[26] , \u_div/QInv[25] ,
         \u_div/QInv[24] , \u_div/QInv[23] , \u_div/QInv[22] ,
         \u_div/QInv[21] , \u_div/QInv[20] , \u_div/QInv[19] ,
         \u_div/QInv[18] , \u_div/QInv[17] , \u_div/QInv[16] ,
         \u_div/QInv[15] , \u_div/QInv[14] , \u_div/QInv[13] ,
         \u_div/QInv[12] , \u_div/QInv[11] , \u_div/QInv[10] , \u_div/QInv[9] ,
         \u_div/QInv[8] , \u_div/QInv[7] , \u_div/QInv[6] , \u_div/QInv[5] ,
         \u_div/QInv[4] , \u_div/QInv[3] , \u_div/QInv[2] , \u_div/QInv[1] ,
         \u_div/QInv[0] , \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] ,
         \u_div/SumTmp[1][3] , \u_div/SumTmp[1][4] , \u_div/SumTmp[2][1] ,
         \u_div/SumTmp[2][2] , \u_div/SumTmp[2][3] , \u_div/SumTmp[2][4] ,
         \u_div/SumTmp[3][1] , \u_div/SumTmp[3][2] , \u_div/SumTmp[3][3] ,
         \u_div/SumTmp[3][4] , \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] ,
         \u_div/SumTmp[4][3] , \u_div/SumTmp[4][4] , \u_div/SumTmp[5][1] ,
         \u_div/SumTmp[5][2] , \u_div/SumTmp[5][3] , \u_div/SumTmp[5][4] ,
         \u_div/SumTmp[6][1] , \u_div/SumTmp[6][2] , \u_div/SumTmp[6][3] ,
         \u_div/SumTmp[6][4] , \u_div/SumTmp[7][1] , \u_div/SumTmp[7][2] ,
         \u_div/SumTmp[7][3] , \u_div/SumTmp[7][4] , \u_div/SumTmp[8][1] ,
         \u_div/SumTmp[8][2] , \u_div/SumTmp[8][3] , \u_div/SumTmp[8][4] ,
         \u_div/SumTmp[9][1] , \u_div/SumTmp[9][2] , \u_div/SumTmp[9][3] ,
         \u_div/SumTmp[9][4] , \u_div/SumTmp[10][1] , \u_div/SumTmp[10][2] ,
         \u_div/SumTmp[10][3] , \u_div/SumTmp[10][4] , \u_div/SumTmp[11][1] ,
         \u_div/SumTmp[11][2] , \u_div/SumTmp[11][3] , \u_div/SumTmp[11][4] ,
         \u_div/SumTmp[12][1] , \u_div/SumTmp[12][2] , \u_div/SumTmp[12][3] ,
         \u_div/SumTmp[12][4] , \u_div/SumTmp[13][1] , \u_div/SumTmp[13][2] ,
         \u_div/SumTmp[13][3] , \u_div/SumTmp[13][4] , \u_div/SumTmp[14][1] ,
         \u_div/SumTmp[14][2] , \u_div/SumTmp[14][3] , \u_div/SumTmp[14][4] ,
         \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] , \u_div/SumTmp[15][3] ,
         \u_div/SumTmp[15][4] , \u_div/SumTmp[16][1] , \u_div/SumTmp[16][2] ,
         \u_div/SumTmp[16][3] , \u_div/SumTmp[16][4] , \u_div/SumTmp[17][1] ,
         \u_div/SumTmp[17][2] , \u_div/SumTmp[17][3] , \u_div/SumTmp[17][4] ,
         \u_div/SumTmp[18][1] , \u_div/SumTmp[18][2] , \u_div/SumTmp[18][3] ,
         \u_div/SumTmp[18][4] , \u_div/SumTmp[19][1] , \u_div/SumTmp[19][2] ,
         \u_div/SumTmp[19][3] , \u_div/SumTmp[19][4] , \u_div/SumTmp[20][1] ,
         \u_div/SumTmp[20][2] , \u_div/SumTmp[20][3] , \u_div/SumTmp[20][4] ,
         \u_div/SumTmp[21][1] , \u_div/SumTmp[21][2] , \u_div/SumTmp[21][3] ,
         \u_div/SumTmp[21][4] , \u_div/SumTmp[22][1] , \u_div/SumTmp[22][2] ,
         \u_div/SumTmp[22][3] , \u_div/SumTmp[22][4] , \u_div/SumTmp[23][1] ,
         \u_div/SumTmp[23][2] , \u_div/SumTmp[23][3] , \u_div/SumTmp[23][4] ,
         \u_div/SumTmp[24][1] , \u_div/SumTmp[24][2] , \u_div/SumTmp[24][3] ,
         \u_div/SumTmp[24][4] , \u_div/SumTmp[25][1] , \u_div/SumTmp[25][2] ,
         \u_div/SumTmp[25][3] , \u_div/SumTmp[25][4] , \u_div/SumTmp[26][1] ,
         \u_div/SumTmp[26][2] , \u_div/SumTmp[26][3] , \u_div/SumTmp[26][4] ,
         \u_div/SumTmp[27][1] , \u_div/SumTmp[27][2] , \u_div/SumTmp[27][3] ,
         \u_div/SumTmp[27][4] , \u_div/SumTmp[28][1] , \u_div/SumTmp[28][2] ,
         \u_div/SumTmp[28][3] , \u_div/SumTmp[28][4] , \u_div/SumTmp[29][1] ,
         \u_div/SumTmp[29][2] , \u_div/SumTmp[29][3] , \u_div/SumTmp[29][4] ,
         \u_div/SumTmp[30][1] , \u_div/SumTmp[30][2] , \u_div/SumTmp[30][3] ,
         \u_div/SumTmp[30][4] , \u_div/SumTmp[31][1] , \u_div/SumTmp[31][2] ,
         \u_div/SumTmp[31][3] , \u_div/SumTmp[31][4] , \u_div/SumTmp[32][1] ,
         \u_div/SumTmp[32][2] , \u_div/SumTmp[32][3] , \u_div/SumTmp[32][4] ,
         \u_div/SumTmp[33][1] , \u_div/SumTmp[33][2] , \u_div/SumTmp[33][3] ,
         \u_div/SumTmp[33][4] , \u_div/SumTmp[34][1] , \u_div/SumTmp[34][2] ,
         \u_div/SumTmp[34][3] , \u_div/SumTmp[34][4] , \u_div/SumTmp[35][1] ,
         \u_div/SumTmp[35][2] , \u_div/SumTmp[35][3] , \u_div/SumTmp[35][4] ,
         \u_div/SumTmp[36][1] , \u_div/SumTmp[36][2] , \u_div/SumTmp[36][3] ,
         \u_div/SumTmp[36][4] , \u_div/SumTmp[37][1] , \u_div/SumTmp[37][2] ,
         \u_div/SumTmp[37][3] , \u_div/SumTmp[37][4] , \u_div/SumTmp[38][1] ,
         \u_div/SumTmp[38][2] , \u_div/SumTmp[38][3] , \u_div/SumTmp[38][4] ,
         \u_div/SumTmp[39][1] , \u_div/SumTmp[39][2] , \u_div/SumTmp[39][3] ,
         \u_div/SumTmp[39][4] , \u_div/SumTmp[40][1] , \u_div/SumTmp[40][2] ,
         \u_div/SumTmp[40][3] , \u_div/SumTmp[40][4] , \u_div/SumTmp[41][1] ,
         \u_div/SumTmp[41][2] , \u_div/SumTmp[41][3] , \u_div/SumTmp[41][4] ,
         \u_div/SumTmp[42][1] , \u_div/SumTmp[42][2] , \u_div/SumTmp[42][3] ,
         \u_div/SumTmp[42][4] , \u_div/SumTmp[43][1] , \u_div/SumTmp[43][2] ,
         \u_div/SumTmp[43][3] , \u_div/SumTmp[43][4] , \u_div/SumTmp[44][1] ,
         \u_div/SumTmp[44][2] , \u_div/SumTmp[44][3] , \u_div/SumTmp[44][4] ,
         \u_div/SumTmp[45][1] , \u_div/SumTmp[45][2] , \u_div/SumTmp[45][3] ,
         \u_div/SumTmp[45][4] , \u_div/SumTmp[46][1] , \u_div/SumTmp[46][2] ,
         \u_div/SumTmp[46][3] , \u_div/SumTmp[46][4] , \u_div/SumTmp[47][1] ,
         \u_div/SumTmp[47][2] , \u_div/SumTmp[47][3] , \u_div/SumTmp[47][4] ,
         \u_div/SumTmp[48][1] , \u_div/SumTmp[48][2] , \u_div/SumTmp[48][3] ,
         \u_div/SumTmp[48][4] , \u_div/SumTmp[49][1] , \u_div/SumTmp[49][2] ,
         \u_div/SumTmp[49][3] , \u_div/SumTmp[49][4] , \u_div/SumTmp[50][1] ,
         \u_div/SumTmp[50][2] , \u_div/SumTmp[50][3] , \u_div/SumTmp[50][4] ,
         \u_div/SumTmp[51][1] , \u_div/SumTmp[51][2] , \u_div/SumTmp[51][3] ,
         \u_div/SumTmp[51][4] , \u_div/SumTmp[52][1] , \u_div/SumTmp[52][2] ,
         \u_div/SumTmp[52][3] , \u_div/SumTmp[52][4] , \u_div/SumTmp[53][1] ,
         \u_div/SumTmp[53][2] , \u_div/SumTmp[53][3] , \u_div/SumTmp[53][4] ,
         \u_div/SumTmp[54][1] , \u_div/SumTmp[54][2] , \u_div/SumTmp[54][3] ,
         \u_div/SumTmp[54][4] , \u_div/SumTmp[55][1] , \u_div/SumTmp[55][2] ,
         \u_div/SumTmp[55][3] , \u_div/SumTmp[55][4] , \u_div/SumTmp[56][1] ,
         \u_div/SumTmp[56][2] , \u_div/SumTmp[56][3] , \u_div/SumTmp[56][4] ,
         \u_div/SumTmp[57][1] , \u_div/SumTmp[57][2] , \u_div/SumTmp[57][3] ,
         \u_div/SumTmp[57][4] , \u_div/SumTmp[58][1] , \u_div/SumTmp[58][2] ,
         \u_div/SumTmp[58][3] , \u_div/SumTmp[58][4] , \u_div/SumTmp[59][3] ,
         \u_div/SumTmp[59][4] , \u_div/CryTmp[0][6] , \u_div/CryTmp[1][6] ,
         \u_div/CryTmp[2][6] , \u_div/CryTmp[3][6] , \u_div/CryTmp[4][6] ,
         \u_div/CryTmp[5][6] , \u_div/CryTmp[6][6] , \u_div/CryTmp[7][6] ,
         \u_div/CryTmp[8][6] , \u_div/CryTmp[9][6] , \u_div/CryTmp[10][6] ,
         \u_div/CryTmp[11][6] , \u_div/CryTmp[12][6] , \u_div/CryTmp[13][6] ,
         \u_div/CryTmp[14][6] , \u_div/CryTmp[15][6] , \u_div/CryTmp[16][6] ,
         \u_div/CryTmp[17][6] , \u_div/CryTmp[18][6] , \u_div/CryTmp[19][6] ,
         \u_div/CryTmp[20][6] , \u_div/CryTmp[21][6] , \u_div/CryTmp[22][6] ,
         \u_div/CryTmp[23][6] , \u_div/CryTmp[24][6] , \u_div/CryTmp[25][6] ,
         \u_div/CryTmp[26][6] , \u_div/CryTmp[27][6] , \u_div/CryTmp[28][6] ,
         \u_div/CryTmp[29][6] , \u_div/CryTmp[30][6] , \u_div/CryTmp[31][6] ,
         \u_div/CryTmp[32][6] , \u_div/CryTmp[33][6] , \u_div/CryTmp[34][6] ,
         \u_div/CryTmp[35][6] , \u_div/CryTmp[36][6] , \u_div/CryTmp[37][6] ,
         \u_div/CryTmp[38][6] , \u_div/CryTmp[39][6] , \u_div/CryTmp[40][6] ,
         \u_div/CryTmp[41][6] , \u_div/CryTmp[42][6] , \u_div/CryTmp[43][6] ,
         \u_div/CryTmp[44][6] , \u_div/CryTmp[45][6] , \u_div/CryTmp[46][6] ,
         \u_div/CryTmp[47][6] , \u_div/CryTmp[48][6] , \u_div/CryTmp[49][6] ,
         \u_div/CryTmp[50][6] , \u_div/CryTmp[51][6] , \u_div/CryTmp[52][6] ,
         \u_div/CryTmp[53][6] , \u_div/CryTmp[54][6] , \u_div/CryTmp[55][6] ,
         \u_div/CryTmp[56][6] , \u_div/CryTmp[57][6] , \u_div/CryTmp[58][6] ,
         \u_div/CryTmp[59][6] , \u_div/PartRem[1][3] , \u_div/PartRem[1][4] ,
         \u_div/PartRem[1][5] , \u_div/PartRem[2][2] , \u_div/PartRem[2][3] ,
         \u_div/PartRem[2][4] , \u_div/PartRem[2][5] , \u_div/PartRem[3][0] ,
         \u_div/PartRem[3][2] , \u_div/PartRem[3][3] , \u_div/PartRem[3][4] ,
         \u_div/PartRem[3][5] , \u_div/PartRem[4][0] , \u_div/PartRem[4][2] ,
         \u_div/PartRem[4][3] , \u_div/PartRem[4][4] , \u_div/PartRem[4][5] ,
         \u_div/PartRem[5][0] , \u_div/PartRem[5][2] , \u_div/PartRem[5][3] ,
         \u_div/PartRem[5][4] , \u_div/PartRem[5][5] , \u_div/PartRem[6][0] ,
         \u_div/PartRem[6][2] , \u_div/PartRem[6][3] , \u_div/PartRem[6][4] ,
         \u_div/PartRem[6][5] , \u_div/PartRem[7][0] , \u_div/PartRem[7][2] ,
         \u_div/PartRem[7][3] , \u_div/PartRem[7][4] , \u_div/PartRem[7][5] ,
         \u_div/PartRem[8][0] , \u_div/PartRem[8][2] , \u_div/PartRem[8][3] ,
         \u_div/PartRem[8][4] , \u_div/PartRem[8][5] , \u_div/PartRem[9][0] ,
         \u_div/PartRem[9][2] , \u_div/PartRem[9][3] , \u_div/PartRem[9][4] ,
         \u_div/PartRem[9][5] , \u_div/PartRem[10][0] , \u_div/PartRem[10][2] ,
         \u_div/PartRem[10][3] , \u_div/PartRem[10][4] ,
         \u_div/PartRem[10][5] , \u_div/PartRem[11][0] ,
         \u_div/PartRem[11][2] , \u_div/PartRem[11][3] ,
         \u_div/PartRem[11][4] , \u_div/PartRem[11][5] ,
         \u_div/PartRem[12][0] , \u_div/PartRem[12][2] ,
         \u_div/PartRem[12][3] , \u_div/PartRem[12][4] ,
         \u_div/PartRem[12][5] , \u_div/PartRem[13][0] ,
         \u_div/PartRem[13][2] , \u_div/PartRem[13][3] ,
         \u_div/PartRem[13][4] , \u_div/PartRem[13][5] ,
         \u_div/PartRem[14][0] , \u_div/PartRem[14][2] ,
         \u_div/PartRem[14][3] , \u_div/PartRem[14][4] ,
         \u_div/PartRem[14][5] , \u_div/PartRem[15][0] ,
         \u_div/PartRem[15][2] , \u_div/PartRem[15][3] ,
         \u_div/PartRem[15][4] , \u_div/PartRem[15][5] ,
         \u_div/PartRem[16][0] , \u_div/PartRem[16][2] ,
         \u_div/PartRem[16][3] , \u_div/PartRem[16][4] ,
         \u_div/PartRem[16][5] , \u_div/PartRem[17][0] ,
         \u_div/PartRem[17][2] , \u_div/PartRem[17][3] ,
         \u_div/PartRem[17][4] , \u_div/PartRem[17][5] ,
         \u_div/PartRem[18][0] , \u_div/PartRem[18][2] ,
         \u_div/PartRem[18][3] , \u_div/PartRem[18][4] ,
         \u_div/PartRem[18][5] , \u_div/PartRem[19][0] ,
         \u_div/PartRem[19][2] , \u_div/PartRem[19][3] ,
         \u_div/PartRem[19][4] , \u_div/PartRem[19][5] ,
         \u_div/PartRem[20][0] , \u_div/PartRem[20][2] ,
         \u_div/PartRem[20][3] , \u_div/PartRem[20][4] ,
         \u_div/PartRem[20][5] , \u_div/PartRem[21][0] ,
         \u_div/PartRem[21][2] , \u_div/PartRem[21][3] ,
         \u_div/PartRem[21][4] , \u_div/PartRem[21][5] ,
         \u_div/PartRem[22][0] , \u_div/PartRem[22][2] ,
         \u_div/PartRem[22][3] , \u_div/PartRem[22][4] ,
         \u_div/PartRem[22][5] , \u_div/PartRem[23][0] ,
         \u_div/PartRem[23][2] , \u_div/PartRem[23][3] ,
         \u_div/PartRem[23][4] , \u_div/PartRem[23][5] ,
         \u_div/PartRem[24][0] , \u_div/PartRem[24][2] ,
         \u_div/PartRem[24][3] , \u_div/PartRem[24][4] ,
         \u_div/PartRem[24][5] , \u_div/PartRem[25][0] ,
         \u_div/PartRem[25][2] , \u_div/PartRem[25][3] ,
         \u_div/PartRem[25][4] , \u_div/PartRem[25][5] ,
         \u_div/PartRem[26][0] , \u_div/PartRem[26][2] ,
         \u_div/PartRem[26][3] , \u_div/PartRem[26][4] ,
         \u_div/PartRem[26][5] , \u_div/PartRem[27][0] ,
         \u_div/PartRem[27][2] , \u_div/PartRem[27][3] ,
         \u_div/PartRem[27][4] , \u_div/PartRem[27][5] ,
         \u_div/PartRem[28][0] , \u_div/PartRem[28][2] ,
         \u_div/PartRem[28][3] , \u_div/PartRem[28][4] ,
         \u_div/PartRem[28][5] , \u_div/PartRem[29][0] ,
         \u_div/PartRem[29][2] , \u_div/PartRem[29][3] ,
         \u_div/PartRem[29][4] , \u_div/PartRem[29][5] ,
         \u_div/PartRem[30][0] , \u_div/PartRem[30][2] ,
         \u_div/PartRem[30][3] , \u_div/PartRem[30][4] ,
         \u_div/PartRem[30][5] , \u_div/PartRem[31][0] ,
         \u_div/PartRem[31][2] , \u_div/PartRem[31][3] ,
         \u_div/PartRem[31][4] , \u_div/PartRem[31][5] ,
         \u_div/PartRem[32][0] , \u_div/PartRem[32][2] ,
         \u_div/PartRem[32][3] , \u_div/PartRem[32][4] ,
         \u_div/PartRem[32][5] , \u_div/PartRem[33][0] ,
         \u_div/PartRem[33][2] , \u_div/PartRem[33][3] ,
         \u_div/PartRem[33][4] , \u_div/PartRem[33][5] ,
         \u_div/PartRem[34][0] , \u_div/PartRem[34][2] ,
         \u_div/PartRem[34][3] , \u_div/PartRem[34][4] ,
         \u_div/PartRem[34][5] , \u_div/PartRem[35][0] ,
         \u_div/PartRem[35][2] , \u_div/PartRem[35][3] ,
         \u_div/PartRem[35][4] , \u_div/PartRem[35][5] ,
         \u_div/PartRem[36][0] , \u_div/PartRem[36][2] ,
         \u_div/PartRem[36][3] , \u_div/PartRem[36][4] ,
         \u_div/PartRem[36][5] , \u_div/PartRem[37][0] ,
         \u_div/PartRem[37][2] , \u_div/PartRem[37][3] ,
         \u_div/PartRem[37][4] , \u_div/PartRem[37][5] ,
         \u_div/PartRem[38][0] , \u_div/PartRem[38][2] ,
         \u_div/PartRem[38][3] , \u_div/PartRem[38][4] ,
         \u_div/PartRem[38][5] , \u_div/PartRem[39][0] ,
         \u_div/PartRem[39][2] , \u_div/PartRem[39][3] ,
         \u_div/PartRem[39][4] , \u_div/PartRem[39][5] ,
         \u_div/PartRem[40][0] , \u_div/PartRem[40][2] ,
         \u_div/PartRem[40][3] , \u_div/PartRem[40][4] ,
         \u_div/PartRem[40][5] , \u_div/PartRem[41][0] ,
         \u_div/PartRem[41][2] , \u_div/PartRem[41][3] ,
         \u_div/PartRem[41][4] , \u_div/PartRem[41][5] ,
         \u_div/PartRem[42][0] , \u_div/PartRem[42][2] ,
         \u_div/PartRem[42][3] , \u_div/PartRem[42][4] ,
         \u_div/PartRem[42][5] , \u_div/PartRem[43][0] ,
         \u_div/PartRem[43][2] , \u_div/PartRem[43][3] ,
         \u_div/PartRem[43][4] , \u_div/PartRem[43][5] ,
         \u_div/PartRem[44][0] , \u_div/PartRem[44][2] ,
         \u_div/PartRem[44][3] , \u_div/PartRem[44][4] ,
         \u_div/PartRem[44][5] , \u_div/PartRem[45][0] ,
         \u_div/PartRem[45][2] , \u_div/PartRem[45][3] ,
         \u_div/PartRem[45][4] , \u_div/PartRem[45][5] ,
         \u_div/PartRem[46][0] , \u_div/PartRem[46][2] ,
         \u_div/PartRem[46][3] , \u_div/PartRem[46][4] ,
         \u_div/PartRem[46][5] , \u_div/PartRem[47][0] ,
         \u_div/PartRem[47][2] , \u_div/PartRem[47][3] ,
         \u_div/PartRem[47][4] , \u_div/PartRem[47][5] ,
         \u_div/PartRem[48][0] , \u_div/PartRem[48][2] ,
         \u_div/PartRem[48][3] , \u_div/PartRem[48][4] ,
         \u_div/PartRem[48][5] , \u_div/PartRem[49][0] ,
         \u_div/PartRem[49][2] , \u_div/PartRem[49][3] ,
         \u_div/PartRem[49][4] , \u_div/PartRem[49][5] ,
         \u_div/PartRem[50][0] , \u_div/PartRem[50][2] ,
         \u_div/PartRem[50][3] , \u_div/PartRem[50][4] ,
         \u_div/PartRem[50][5] , \u_div/PartRem[51][0] ,
         \u_div/PartRem[51][2] , \u_div/PartRem[51][3] ,
         \u_div/PartRem[51][4] , \u_div/PartRem[51][5] ,
         \u_div/PartRem[52][0] , \u_div/PartRem[52][2] ,
         \u_div/PartRem[52][3] , \u_div/PartRem[52][4] ,
         \u_div/PartRem[52][5] , \u_div/PartRem[53][0] ,
         \u_div/PartRem[53][2] , \u_div/PartRem[53][3] ,
         \u_div/PartRem[53][4] , \u_div/PartRem[53][5] ,
         \u_div/PartRem[54][0] , \u_div/PartRem[54][2] ,
         \u_div/PartRem[54][3] , \u_div/PartRem[54][4] ,
         \u_div/PartRem[54][5] , \u_div/PartRem[55][0] ,
         \u_div/PartRem[55][2] , \u_div/PartRem[55][3] ,
         \u_div/PartRem[55][4] , \u_div/PartRem[55][5] ,
         \u_div/PartRem[56][0] , \u_div/PartRem[56][2] ,
         \u_div/PartRem[56][3] , \u_div/PartRem[56][4] ,
         \u_div/PartRem[56][5] , \u_div/PartRem[57][0] ,
         \u_div/PartRem[57][2] , \u_div/PartRem[57][3] ,
         \u_div/PartRem[57][4] , \u_div/PartRem[57][5] ,
         \u_div/PartRem[58][0] , \u_div/PartRem[58][2] ,
         \u_div/PartRem[58][3] , \u_div/PartRem[58][4] ,
         \u_div/PartRem[58][5] , \u_div/PartRem[59][0] ,
         \u_div/PartRem[59][2] , \u_div/PartRem[59][3] ,
         \u_div/PartRem[59][4] , \u_div/PartRem[59][5] ,
         \u_div/PartRem[60][0] , \u_div/PartRem[61][0] ,
         \u_div/PartRem[62][0] , \u_div/PartRem[63][0] ,
         \u_div/PartRem[64][0] , \u_div/u_add_PartRem_2_1/n3 ,
         \u_div/u_add_PartRem_2_1/n2 , \u_div/u_add_PartRem_2_2/n3 ,
         \u_div/u_add_PartRem_2_2/n2 , \u_div/u_add_PartRem_2_3/n3 ,
         \u_div/u_add_PartRem_2_3/n2 , \u_div/u_add_PartRem_2_4/n3 ,
         \u_div/u_add_PartRem_2_4/n2 , \u_div/u_add_PartRem_2_5/n3 ,
         \u_div/u_add_PartRem_2_5/n2 , \u_div/u_add_PartRem_2_6/n3 ,
         \u_div/u_add_PartRem_2_6/n2 , \u_div/u_add_PartRem_2_7/n3 ,
         \u_div/u_add_PartRem_2_7/n2 , \u_div/u_add_PartRem_2_8/n3 ,
         \u_div/u_add_PartRem_2_8/n2 , \u_div/u_add_PartRem_2_9/n3 ,
         \u_div/u_add_PartRem_2_9/n2 , \u_div/u_add_PartRem_2_10/n3 ,
         \u_div/u_add_PartRem_2_10/n2 , \u_div/u_add_PartRem_2_11/n3 ,
         \u_div/u_add_PartRem_2_11/n2 , \u_div/u_add_PartRem_2_12/n3 ,
         \u_div/u_add_PartRem_2_12/n2 , \u_div/u_add_PartRem_2_13/n3 ,
         \u_div/u_add_PartRem_2_13/n2 , \u_div/u_add_PartRem_2_14/n3 ,
         \u_div/u_add_PartRem_2_14/n2 , \u_div/u_add_PartRem_2_15/n3 ,
         \u_div/u_add_PartRem_2_15/n2 , \u_div/u_add_PartRem_2_16/n3 ,
         \u_div/u_add_PartRem_2_16/n2 , \u_div/u_add_PartRem_2_17/n3 ,
         \u_div/u_add_PartRem_2_17/n2 , \u_div/u_add_PartRem_2_18/n3 ,
         \u_div/u_add_PartRem_2_18/n2 , \u_div/u_add_PartRem_2_19/n3 ,
         \u_div/u_add_PartRem_2_19/n2 , \u_div/u_add_PartRem_2_20/n3 ,
         \u_div/u_add_PartRem_2_20/n2 , \u_div/u_add_PartRem_2_21/n3 ,
         \u_div/u_add_PartRem_2_21/n2 , \u_div/u_add_PartRem_2_22/n3 ,
         \u_div/u_add_PartRem_2_22/n2 , \u_div/u_add_PartRem_2_23/n3 ,
         \u_div/u_add_PartRem_2_23/n2 , \u_div/u_add_PartRem_2_24/n3 ,
         \u_div/u_add_PartRem_2_24/n2 , \u_div/u_add_PartRem_2_25/n3 ,
         \u_div/u_add_PartRem_2_25/n2 , \u_div/u_add_PartRem_2_26/n3 ,
         \u_div/u_add_PartRem_2_26/n2 , \u_div/u_add_PartRem_2_27/n3 ,
         \u_div/u_add_PartRem_2_27/n2 , \u_div/u_add_PartRem_2_28/n3 ,
         \u_div/u_add_PartRem_2_28/n2 , \u_div/u_add_PartRem_2_29/n3 ,
         \u_div/u_add_PartRem_2_29/n2 , \u_div/u_add_PartRem_2_30/n3 ,
         \u_div/u_add_PartRem_2_30/n2 , \u_div/u_add_PartRem_2_31/n3 ,
         \u_div/u_add_PartRem_2_31/n2 , \u_div/u_add_PartRem_2_32/n3 ,
         \u_div/u_add_PartRem_2_32/n2 , \u_div/u_add_PartRem_2_33/n3 ,
         \u_div/u_add_PartRem_2_33/n2 , \u_div/u_add_PartRem_2_34/n3 ,
         \u_div/u_add_PartRem_2_34/n2 , \u_div/u_add_PartRem_2_35/n3 ,
         \u_div/u_add_PartRem_2_35/n2 , \u_div/u_add_PartRem_2_36/n3 ,
         \u_div/u_add_PartRem_2_36/n2 , \u_div/u_add_PartRem_2_37/n3 ,
         \u_div/u_add_PartRem_2_37/n2 , \u_div/u_add_PartRem_2_38/n3 ,
         \u_div/u_add_PartRem_2_38/n2 , \u_div/u_add_PartRem_2_39/n3 ,
         \u_div/u_add_PartRem_2_39/n2 , \u_div/u_add_PartRem_2_40/n3 ,
         \u_div/u_add_PartRem_2_40/n2 , \u_div/u_add_PartRem_2_41/n3 ,
         \u_div/u_add_PartRem_2_41/n2 , \u_div/u_add_PartRem_2_42/n3 ,
         \u_div/u_add_PartRem_2_42/n2 , \u_div/u_add_PartRem_2_43/n3 ,
         \u_div/u_add_PartRem_2_43/n2 , \u_div/u_add_PartRem_2_44/n3 ,
         \u_div/u_add_PartRem_2_44/n2 , \u_div/u_add_PartRem_2_45/n3 ,
         \u_div/u_add_PartRem_2_45/n2 , \u_div/u_add_PartRem_2_46/n3 ,
         \u_div/u_add_PartRem_2_46/n2 , \u_div/u_add_PartRem_2_47/n3 ,
         \u_div/u_add_PartRem_2_47/n2 , \u_div/u_add_PartRem_2_48/n3 ,
         \u_div/u_add_PartRem_2_48/n2 , \u_div/u_add_PartRem_2_49/n3 ,
         \u_div/u_add_PartRem_2_49/n2 , \u_div/u_add_PartRem_2_50/n3 ,
         \u_div/u_add_PartRem_2_50/n2 , \u_div/u_add_PartRem_2_51/n3 ,
         \u_div/u_add_PartRem_2_51/n2 , \u_div/u_add_PartRem_2_52/n3 ,
         \u_div/u_add_PartRem_2_52/n2 , \u_div/u_add_PartRem_2_53/n3 ,
         \u_div/u_add_PartRem_2_53/n2 , \u_div/u_add_PartRem_2_54/n3 ,
         \u_div/u_add_PartRem_2_54/n2 , \u_div/u_add_PartRem_2_55/n3 ,
         \u_div/u_add_PartRem_2_55/n2 , \u_div/u_add_PartRem_2_56/n3 ,
         \u_div/u_add_PartRem_2_56/n2 , \u_div/u_add_PartRem_2_57/n3 ,
         \u_div/u_add_PartRem_2_57/n2 , \u_div/u_add_PartRem_2_58/n3 ,
         \u_div/u_add_PartRem_2_58/n2 , n1, n2, n3, n4, n5, n6, n7, n8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign \u_div/QInv[63]  = a[63];

  GSIM_DW01_absval_1 \u_div/u_absval_AAbs  ( .A({n3, a[62:0]}), .ABSVAL({
        \u_div/PartRem[64][0] , \u_div/PartRem[63][0] , \u_div/PartRem[62][0] , 
        \u_div/PartRem[61][0] , \u_div/PartRem[60][0] , \u_div/PartRem[59][0] , 
        \u_div/PartRem[58][0] , \u_div/PartRem[57][0] , \u_div/PartRem[56][0] , 
        \u_div/PartRem[55][0] , \u_div/PartRem[54][0] , \u_div/PartRem[53][0] , 
        \u_div/PartRem[52][0] , \u_div/PartRem[51][0] , \u_div/PartRem[50][0] , 
        \u_div/PartRem[49][0] , \u_div/PartRem[48][0] , \u_div/PartRem[47][0] , 
        \u_div/PartRem[46][0] , \u_div/PartRem[45][0] , \u_div/PartRem[44][0] , 
        \u_div/PartRem[43][0] , \u_div/PartRem[42][0] , \u_div/PartRem[41][0] , 
        \u_div/PartRem[40][0] , \u_div/PartRem[39][0] , \u_div/PartRem[38][0] , 
        \u_div/PartRem[37][0] , \u_div/PartRem[36][0] , \u_div/PartRem[35][0] , 
        \u_div/PartRem[34][0] , \u_div/PartRem[33][0] , \u_div/PartRem[32][0] , 
        \u_div/PartRem[31][0] , \u_div/PartRem[30][0] , \u_div/PartRem[29][0] , 
        \u_div/PartRem[28][0] , \u_div/PartRem[27][0] , \u_div/PartRem[26][0] , 
        \u_div/PartRem[25][0] , \u_div/PartRem[24][0] , \u_div/PartRem[23][0] , 
        \u_div/PartRem[22][0] , \u_div/PartRem[21][0] , \u_div/PartRem[20][0] , 
        \u_div/PartRem[19][0] , \u_div/PartRem[18][0] , \u_div/PartRem[17][0] , 
        \u_div/PartRem[16][0] , \u_div/PartRem[15][0] , \u_div/PartRem[14][0] , 
        \u_div/PartRem[13][0] , \u_div/PartRem[12][0] , \u_div/PartRem[11][0] , 
        \u_div/PartRem[10][0] , \u_div/PartRem[9][0] , \u_div/PartRem[8][0] , 
        \u_div/PartRem[7][0] , \u_div/PartRem[6][0] , \u_div/PartRem[5][0] , 
        \u_div/PartRem[4][0] , \u_div/PartRem[3][0] , SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1}) );
  GSIM_DW_inc_1 \u_div/u_inc_QInc  ( .carry_in(n5), .a({n3, n3, n3, n4, 
        \u_div/QInv[59] , \u_div/QInv[58] , \u_div/QInv[57] , \u_div/QInv[56] , 
        \u_div/QInv[55] , \u_div/QInv[54] , \u_div/QInv[53] , \u_div/QInv[52] , 
        \u_div/QInv[51] , \u_div/QInv[50] , \u_div/QInv[49] , \u_div/QInv[48] , 
        \u_div/QInv[47] , \u_div/QInv[46] , \u_div/QInv[45] , \u_div/QInv[44] , 
        \u_div/QInv[43] , \u_div/QInv[42] , \u_div/QInv[41] , \u_div/QInv[40] , 
        \u_div/QInv[39] , \u_div/QInv[38] , \u_div/QInv[37] , \u_div/QInv[36] , 
        \u_div/QInv[35] , \u_div/QInv[34] , \u_div/QInv[33] , \u_div/QInv[32] , 
        \u_div/QInv[31] , \u_div/QInv[30] , \u_div/QInv[29] , \u_div/QInv[28] , 
        \u_div/QInv[27] , \u_div/QInv[26] , \u_div/QInv[25] , \u_div/QInv[24] , 
        \u_div/QInv[23] , \u_div/QInv[22] , \u_div/QInv[21] , \u_div/QInv[20] , 
        \u_div/QInv[19] , \u_div/QInv[18] , \u_div/QInv[17] , \u_div/QInv[16] , 
        \u_div/QInv[15] , \u_div/QInv[14] , \u_div/QInv[13] , \u_div/QInv[12] , 
        \u_div/QInv[11] , \u_div/QInv[10] , \u_div/QInv[9] , \u_div/QInv[8] , 
        \u_div/QInv[7] , \u_div/QInv[6] , \u_div/QInv[5] , \u_div/QInv[4] , 
        \u_div/QInv[3] , \u_div/QInv[2] , \u_div/QInv[1] , \u_div/QInv[0] }), 
        .sum(quotient) );
  ADDHXL \u_div/u_add_PartRem_2_3/U3  ( .A(\u_div/PartRem[4][4] ), .B(
        \u_div/u_add_PartRem_2_3/n3 ), .CO(\u_div/u_add_PartRem_2_3/n2 ), .S(
        \u_div/SumTmp[3][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_12/U3  ( .A(\u_div/PartRem[13][4] ), .B(
        \u_div/u_add_PartRem_2_12/n3 ), .CO(\u_div/u_add_PartRem_2_12/n2 ), 
        .S(\u_div/SumTmp[12][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_17/U3  ( .A(\u_div/PartRem[18][4] ), .B(
        \u_div/u_add_PartRem_2_17/n3 ), .CO(\u_div/u_add_PartRem_2_17/n2 ), 
        .S(\u_div/SumTmp[17][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_22/U3  ( .A(\u_div/PartRem[23][4] ), .B(
        \u_div/u_add_PartRem_2_22/n3 ), .CO(\u_div/u_add_PartRem_2_22/n2 ), 
        .S(\u_div/SumTmp[22][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_27/U3  ( .A(\u_div/PartRem[28][4] ), .B(
        \u_div/u_add_PartRem_2_27/n3 ), .CO(\u_div/u_add_PartRem_2_27/n2 ), 
        .S(\u_div/SumTmp[27][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_32/U3  ( .A(\u_div/PartRem[33][4] ), .B(
        \u_div/u_add_PartRem_2_32/n3 ), .CO(\u_div/u_add_PartRem_2_32/n2 ), 
        .S(\u_div/SumTmp[32][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_37/U3  ( .A(\u_div/PartRem[38][4] ), .B(
        \u_div/u_add_PartRem_2_37/n3 ), .CO(\u_div/u_add_PartRem_2_37/n2 ), 
        .S(\u_div/SumTmp[37][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_42/U3  ( .A(\u_div/PartRem[43][4] ), .B(
        \u_div/u_add_PartRem_2_42/n3 ), .CO(\u_div/u_add_PartRem_2_42/n2 ), 
        .S(\u_div/SumTmp[42][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_47/U3  ( .A(\u_div/PartRem[48][4] ), .B(
        \u_div/u_add_PartRem_2_47/n3 ), .CO(\u_div/u_add_PartRem_2_47/n2 ), 
        .S(\u_div/SumTmp[47][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_52/U3  ( .A(\u_div/PartRem[53][4] ), .B(
        \u_div/u_add_PartRem_2_52/n3 ), .CO(\u_div/u_add_PartRem_2_52/n2 ), 
        .S(\u_div/SumTmp[52][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_0  ( .A(\u_div/PartRem[4][0] ), .B(
        \u_div/PartRem[4][0] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/SumTmp[2][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_2_1  ( .A(\u_div/SumTmp[2][1] ), .B(
        \u_div/SumTmp[2][1] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_0  ( .A(\u_div/PartRem[7][0] ), .B(
        \u_div/PartRem[7][0] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/SumTmp[5][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_0  ( .A(\u_div/PartRem[8][0] ), .B(
        \u_div/PartRem[8][0] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/SumTmp[6][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_8_0  ( .A(\u_div/PartRem[9][0] ), .B(
        \u_div/PartRem[9][0] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/SumTmp[7][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_0  ( .A(\u_div/PartRem[11][0] ), .B(
        \u_div/PartRem[11][0] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/SumTmp[9][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_0  ( .A(\u_div/PartRem[12][0] ), .B(
        \u_div/PartRem[12][0] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/SumTmp[10][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_0  ( .A(\u_div/PartRem[13][0] ), .B(
        \u_div/PartRem[13][0] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/SumTmp[11][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_0  ( .A(\u_div/PartRem[14][0] ), .B(
        \u_div/PartRem[14][0] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/SumTmp[12][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_0  ( .A(\u_div/PartRem[16][0] ), .B(
        \u_div/PartRem[16][0] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/SumTmp[14][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_0  ( .A(\u_div/PartRem[17][0] ), .B(
        \u_div/PartRem[17][0] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/SumTmp[15][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_0  ( .A(\u_div/PartRem[18][0] ), .B(
        \u_div/PartRem[18][0] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/SumTmp[16][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_0  ( .A(\u_div/PartRem[19][0] ), .B(
        \u_div/PartRem[19][0] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/SumTmp[17][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_0  ( .A(\u_div/PartRem[21][0] ), .B(
        \u_div/PartRem[21][0] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/SumTmp[19][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_0  ( .A(\u_div/PartRem[22][0] ), .B(
        \u_div/PartRem[22][0] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/SumTmp[20][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_0  ( .A(\u_div/PartRem[23][0] ), .B(
        \u_div/PartRem[23][0] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/SumTmp[21][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_0  ( .A(\u_div/PartRem[24][0] ), .B(
        \u_div/PartRem[24][0] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/SumTmp[22][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_0  ( .A(\u_div/PartRem[26][0] ), .B(
        \u_div/PartRem[26][0] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/SumTmp[24][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_0  ( .A(\u_div/PartRem[27][0] ), .B(
        \u_div/PartRem[27][0] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/SumTmp[25][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_0  ( .A(\u_div/PartRem[28][0] ), .B(
        \u_div/PartRem[28][0] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/SumTmp[26][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_0  ( .A(\u_div/PartRem[29][0] ), .B(
        \u_div/PartRem[29][0] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/SumTmp[27][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_0  ( .A(\u_div/PartRem[31][0] ), .B(
        \u_div/PartRem[31][0] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/SumTmp[29][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_0  ( .A(\u_div/PartRem[32][0] ), .B(
        \u_div/PartRem[32][0] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/SumTmp[30][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_0  ( .A(\u_div/PartRem[33][0] ), .B(
        \u_div/PartRem[33][0] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/SumTmp[31][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_0  ( .A(\u_div/PartRem[34][0] ), .B(
        \u_div/PartRem[34][0] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/SumTmp[32][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_0  ( .A(\u_div/PartRem[36][0] ), .B(
        \u_div/PartRem[36][0] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/SumTmp[34][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_0  ( .A(\u_div/PartRem[37][0] ), .B(
        \u_div/PartRem[37][0] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/SumTmp[35][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_0  ( .A(\u_div/PartRem[38][0] ), .B(
        \u_div/PartRem[38][0] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/SumTmp[36][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_0  ( .A(\u_div/PartRem[39][0] ), .B(
        \u_div/PartRem[39][0] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/SumTmp[37][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_0  ( .A(\u_div/PartRem[41][0] ), .B(
        \u_div/PartRem[41][0] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/SumTmp[39][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_0  ( .A(\u_div/PartRem[42][0] ), .B(
        \u_div/PartRem[42][0] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/SumTmp[40][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_0  ( .A(\u_div/PartRem[43][0] ), .B(
        \u_div/PartRem[43][0] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/SumTmp[41][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_0  ( .A(\u_div/PartRem[44][0] ), .B(
        \u_div/PartRem[44][0] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/SumTmp[42][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_0  ( .A(\u_div/PartRem[46][0] ), .B(
        \u_div/PartRem[46][0] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/SumTmp[44][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_0  ( .A(\u_div/PartRem[47][0] ), .B(
        \u_div/PartRem[47][0] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/SumTmp[45][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_0  ( .A(\u_div/PartRem[48][0] ), .B(
        \u_div/PartRem[48][0] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/SumTmp[46][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_0  ( .A(\u_div/PartRem[49][0] ), .B(
        \u_div/PartRem[49][0] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/SumTmp[47][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_0  ( .A(\u_div/PartRem[51][0] ), .B(
        \u_div/PartRem[51][0] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/SumTmp[49][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_0  ( .A(\u_div/PartRem[52][0] ), .B(
        \u_div/PartRem[52][0] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/SumTmp[50][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_0  ( .A(\u_div/PartRem[53][0] ), .B(
        \u_div/PartRem[53][0] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/SumTmp[51][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_0  ( .A(\u_div/PartRem[54][0] ), .B(
        \u_div/PartRem[54][0] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/SumTmp[52][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_0  ( .A(\u_div/PartRem[56][0] ), .B(
        \u_div/PartRem[56][0] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/SumTmp[54][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_54_1  ( .A(\u_div/SumTmp[54][1] ), .B(
        \u_div/SumTmp[54][1] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_0  ( .A(\u_div/PartRem[57][0] ), .B(
        \u_div/PartRem[57][0] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/SumTmp[55][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_55_1  ( .A(\u_div/SumTmp[55][1] ), .B(
        \u_div/SumTmp[55][1] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_0  ( .A(\u_div/PartRem[58][0] ), .B(
        \u_div/PartRem[58][0] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/SumTmp[56][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_56_1  ( .A(\u_div/SumTmp[56][1] ), .B(
        \u_div/SumTmp[56][1] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_0  ( .A(\u_div/PartRem[59][0] ), .B(
        \u_div/PartRem[59][0] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/SumTmp[57][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_57_1  ( .A(\u_div/SumTmp[57][1] ), .B(
        \u_div/SumTmp[57][1] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_0  ( .A(\u_div/PartRem[60][0] ), .B(
        \u_div/PartRem[60][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/SumTmp[58][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_58_1  ( .A(\u_div/SumTmp[58][1] ), .B(
        \u_div/SumTmp[58][1] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_9_0  ( .A(\u_div/PartRem[10][0] ), .B(
        \u_div/PartRem[10][0] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/SumTmp[8][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_0  ( .A(\u_div/PartRem[15][0] ), .B(
        \u_div/PartRem[15][0] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/SumTmp[13][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_0  ( .A(\u_div/PartRem[20][0] ), .B(
        \u_div/PartRem[20][0] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/SumTmp[18][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_0  ( .A(\u_div/PartRem[25][0] ), .B(
        \u_div/PartRem[25][0] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/SumTmp[23][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_0  ( .A(\u_div/PartRem[30][0] ), .B(
        \u_div/PartRem[30][0] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/SumTmp[28][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_0  ( .A(\u_div/PartRem[35][0] ), .B(
        \u_div/PartRem[35][0] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/SumTmp[33][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_0  ( .A(\u_div/PartRem[40][0] ), .B(
        \u_div/PartRem[40][0] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/SumTmp[38][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_0  ( .A(\u_div/PartRem[45][0] ), .B(
        \u_div/PartRem[45][0] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/SumTmp[43][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_0  ( .A(\u_div/PartRem[50][0] ), .B(
        \u_div/PartRem[50][0] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/SumTmp[48][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_0  ( .A(\u_div/PartRem[55][0] ), .B(
        \u_div/PartRem[55][0] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/SumTmp[53][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_0  ( .A(\u_div/PartRem[6][0] ), .B(
        \u_div/PartRem[6][0] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/SumTmp[4][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_59_1  ( .A(\u_div/PartRem[61][0] ), .B(
        \u_div/PartRem[61][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_0  ( .A(\u_div/PartRem[5][0] ), .B(
        \u_div/PartRem[5][0] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/SumTmp[3][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_3  ( .A(\u_div/PartRem[5][3] ), .B(
        \u_div/SumTmp[4][3] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_3  ( .A(\u_div/PartRem[6][3] ), .B(
        \u_div/SumTmp[5][3] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_3  ( .A(\u_div/PartRem[7][3] ), .B(
        \u_div/SumTmp[6][3] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_3  ( .A(\u_div/PartRem[8][3] ), .B(
        \u_div/SumTmp[7][3] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_8_3  ( .A(\u_div/PartRem[9][3] ), .B(
        \u_div/SumTmp[8][3] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_9_3  ( .A(\u_div/PartRem[10][3] ), .B(
        \u_div/SumTmp[9][3] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_3  ( .A(\u_div/PartRem[11][3] ), .B(
        \u_div/SumTmp[10][3] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_3  ( .A(\u_div/PartRem[12][3] ), .B(
        \u_div/SumTmp[11][3] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_3  ( .A(\u_div/PartRem[13][3] ), .B(
        \u_div/SumTmp[12][3] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_3  ( .A(\u_div/PartRem[14][3] ), .B(
        \u_div/SumTmp[13][3] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_3  ( .A(\u_div/PartRem[15][3] ), .B(
        \u_div/SumTmp[14][3] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_3  ( .A(\u_div/PartRem[16][3] ), .B(
        \u_div/SumTmp[15][3] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_3  ( .A(\u_div/PartRem[17][3] ), .B(
        \u_div/SumTmp[16][3] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_3  ( .A(\u_div/PartRem[18][3] ), .B(
        \u_div/SumTmp[17][3] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_3  ( .A(\u_div/PartRem[19][3] ), .B(
        \u_div/SumTmp[18][3] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_3  ( .A(\u_div/PartRem[20][3] ), .B(
        \u_div/SumTmp[19][3] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_3  ( .A(\u_div/PartRem[21][3] ), .B(
        \u_div/SumTmp[20][3] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_3  ( .A(\u_div/PartRem[22][3] ), .B(
        \u_div/SumTmp[21][3] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_3  ( .A(\u_div/PartRem[23][3] ), .B(
        \u_div/SumTmp[22][3] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_3  ( .A(\u_div/PartRem[24][3] ), .B(
        \u_div/SumTmp[23][3] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_3  ( .A(\u_div/PartRem[25][3] ), .B(
        \u_div/SumTmp[24][3] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_3  ( .A(\u_div/PartRem[26][3] ), .B(
        \u_div/SumTmp[25][3] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_3  ( .A(\u_div/PartRem[27][3] ), .B(
        \u_div/SumTmp[26][3] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_3  ( .A(\u_div/PartRem[28][3] ), .B(
        \u_div/SumTmp[27][3] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_3  ( .A(\u_div/PartRem[29][3] ), .B(
        \u_div/SumTmp[28][3] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_3  ( .A(\u_div/PartRem[30][3] ), .B(
        \u_div/SumTmp[29][3] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_3  ( .A(\u_div/PartRem[31][3] ), .B(
        \u_div/SumTmp[30][3] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_3  ( .A(\u_div/PartRem[32][3] ), .B(
        \u_div/SumTmp[31][3] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_3  ( .A(\u_div/PartRem[33][3] ), .B(
        \u_div/SumTmp[32][3] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_3  ( .A(\u_div/PartRem[34][3] ), .B(
        \u_div/SumTmp[33][3] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_3  ( .A(\u_div/PartRem[35][3] ), .B(
        \u_div/SumTmp[34][3] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_3  ( .A(\u_div/PartRem[36][3] ), .B(
        \u_div/SumTmp[35][3] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_3  ( .A(\u_div/PartRem[37][3] ), .B(
        \u_div/SumTmp[36][3] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_3  ( .A(\u_div/PartRem[38][3] ), .B(
        \u_div/SumTmp[37][3] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_3  ( .A(\u_div/PartRem[39][3] ), .B(
        \u_div/SumTmp[38][3] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_3  ( .A(\u_div/PartRem[40][3] ), .B(
        \u_div/SumTmp[39][3] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_3  ( .A(\u_div/PartRem[41][3] ), .B(
        \u_div/SumTmp[40][3] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_3  ( .A(\u_div/PartRem[42][3] ), .B(
        \u_div/SumTmp[41][3] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_3  ( .A(\u_div/PartRem[43][3] ), .B(
        \u_div/SumTmp[42][3] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_3  ( .A(\u_div/PartRem[44][3] ), .B(
        \u_div/SumTmp[43][3] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_3  ( .A(\u_div/PartRem[45][3] ), .B(
        \u_div/SumTmp[44][3] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_3  ( .A(\u_div/PartRem[46][3] ), .B(
        \u_div/SumTmp[45][3] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_3  ( .A(\u_div/PartRem[47][3] ), .B(
        \u_div/SumTmp[46][3] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_3  ( .A(\u_div/PartRem[48][3] ), .B(
        \u_div/SumTmp[47][3] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_3  ( .A(\u_div/PartRem[49][3] ), .B(
        \u_div/SumTmp[48][3] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_3  ( .A(\u_div/PartRem[50][3] ), .B(
        \u_div/SumTmp[49][3] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_3  ( .A(\u_div/PartRem[51][3] ), .B(
        \u_div/SumTmp[50][3] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_3  ( .A(\u_div/PartRem[52][3] ), .B(
        \u_div/SumTmp[51][3] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_3  ( .A(\u_div/PartRem[53][3] ), .B(
        \u_div/SumTmp[52][3] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_3  ( .A(\u_div/PartRem[54][3] ), .B(
        \u_div/SumTmp[53][3] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_3  ( .A(\u_div/PartRem[55][3] ), .B(
        \u_div/SumTmp[54][3] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_3  ( .A(\u_div/PartRem[56][3] ), .B(
        \u_div/SumTmp[55][3] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_3  ( .A(\u_div/PartRem[57][3] ), .B(
        \u_div/SumTmp[56][3] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_3  ( .A(\u_div/PartRem[58][3] ), .B(
        \u_div/SumTmp[57][3] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_3  ( .A(\u_div/PartRem[59][3] ), .B(
        \u_div/SumTmp[58][3] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_3  ( .A(\u_div/PartRem[63][0] ), .B(
        \u_div/SumTmp[59][3] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_3  ( .A(\u_div/PartRem[4][3] ), .B(
        \u_div/SumTmp[3][3] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_4  ( .A(\u_div/PartRem[64][0] ), .B(
        \u_div/SumTmp[59][4] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_0  ( .A(\u_div/PartRem[3][0] ), .B(
        \u_div/PartRem[3][0] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/SumTmp[1][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_4_1  ( .A(\u_div/SumTmp[4][1] ), .B(
        \u_div/SumTmp[4][1] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_5_1  ( .A(\u_div/SumTmp[5][1] ), .B(
        \u_div/SumTmp[5][1] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_6_1  ( .A(\u_div/SumTmp[6][1] ), .B(
        \u_div/SumTmp[6][1] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_10_1  ( .A(\u_div/SumTmp[10][1] ), .B(
        \u_div/SumTmp[10][1] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_7_1  ( .A(\u_div/SumTmp[7][1] ), .B(
        \u_div/SumTmp[7][1] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_9_1  ( .A(\u_div/SumTmp[9][1] ), .B(
        \u_div/SumTmp[9][1] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_8_1  ( .A(\u_div/SumTmp[8][1] ), .B(
        \u_div/SumTmp[8][1] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_11_1  ( .A(\u_div/SumTmp[11][1] ), .B(
        \u_div/SumTmp[11][1] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_12_1  ( .A(\u_div/SumTmp[12][1] ), .B(
        \u_div/SumTmp[12][1] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_13_1  ( .A(\u_div/SumTmp[13][1] ), .B(
        \u_div/SumTmp[13][1] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_22_1  ( .A(\u_div/SumTmp[22][1] ), .B(
        \u_div/SumTmp[22][1] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_23_1  ( .A(\u_div/SumTmp[23][1] ), .B(
        \u_div/SumTmp[23][1] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_24_1  ( .A(\u_div/SumTmp[24][1] ), .B(
        \u_div/SumTmp[24][1] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_25_1  ( .A(\u_div/SumTmp[25][1] ), .B(
        \u_div/SumTmp[25][1] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_21_1  ( .A(\u_div/SumTmp[21][1] ), .B(
        \u_div/SumTmp[21][1] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_14_1  ( .A(\u_div/SumTmp[14][1] ), .B(
        \u_div/SumTmp[14][1] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_26_1  ( .A(\u_div/SumTmp[26][1] ), .B(
        \u_div/SumTmp[26][1] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_20_1  ( .A(\u_div/SumTmp[20][1] ), .B(
        \u_div/SumTmp[20][1] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_15_1  ( .A(\u_div/SumTmp[15][1] ), .B(
        \u_div/SumTmp[15][1] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_27_1  ( .A(\u_div/SumTmp[27][1] ), .B(
        \u_div/SumTmp[27][1] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_16_1  ( .A(\u_div/SumTmp[16][1] ), .B(
        \u_div/SumTmp[16][1] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_19_1  ( .A(\u_div/SumTmp[19][1] ), .B(
        \u_div/SumTmp[19][1] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_17_1  ( .A(\u_div/SumTmp[17][1] ), .B(
        \u_div/SumTmp[17][1] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_18_1  ( .A(\u_div/SumTmp[18][1] ), .B(
        \u_div/SumTmp[18][1] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_28_1  ( .A(\u_div/SumTmp[28][1] ), .B(
        \u_div/SumTmp[28][1] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_29_1  ( .A(\u_div/SumTmp[29][1] ), .B(
        \u_div/SumTmp[29][1] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_30_1  ( .A(\u_div/SumTmp[30][1] ), .B(
        \u_div/SumTmp[30][1] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_31_1  ( .A(\u_div/SumTmp[31][1] ), .B(
        \u_div/SumTmp[31][1] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_32_1  ( .A(\u_div/SumTmp[32][1] ), .B(
        \u_div/SumTmp[32][1] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_33_1  ( .A(\u_div/SumTmp[33][1] ), .B(
        \u_div/SumTmp[33][1] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_34_1  ( .A(\u_div/SumTmp[34][1] ), .B(
        \u_div/SumTmp[34][1] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_35_1  ( .A(\u_div/SumTmp[35][1] ), .B(
        \u_div/SumTmp[35][1] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_36_1  ( .A(\u_div/SumTmp[36][1] ), .B(
        \u_div/SumTmp[36][1] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_37_1  ( .A(\u_div/SumTmp[37][1] ), .B(
        \u_div/SumTmp[37][1] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_38_1  ( .A(\u_div/SumTmp[38][1] ), .B(
        \u_div/SumTmp[38][1] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_39_1  ( .A(\u_div/SumTmp[39][1] ), .B(
        \u_div/SumTmp[39][1] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_40_1  ( .A(\u_div/SumTmp[40][1] ), .B(
        \u_div/SumTmp[40][1] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_41_1  ( .A(\u_div/SumTmp[41][1] ), .B(
        \u_div/SumTmp[41][1] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_42_1  ( .A(\u_div/SumTmp[42][1] ), .B(
        \u_div/SumTmp[42][1] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_43_1  ( .A(\u_div/SumTmp[43][1] ), .B(
        \u_div/SumTmp[43][1] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_44_1  ( .A(\u_div/SumTmp[44][1] ), .B(
        \u_div/SumTmp[44][1] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_45_1  ( .A(\u_div/SumTmp[45][1] ), .B(
        \u_div/SumTmp[45][1] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_46_1  ( .A(\u_div/SumTmp[46][1] ), .B(
        \u_div/SumTmp[46][1] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_47_1  ( .A(\u_div/SumTmp[47][1] ), .B(
        \u_div/SumTmp[47][1] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_51_1  ( .A(\u_div/SumTmp[51][1] ), .B(
        \u_div/SumTmp[51][1] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_48_1  ( .A(\u_div/SumTmp[48][1] ), .B(
        \u_div/SumTmp[48][1] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_49_1  ( .A(\u_div/SumTmp[49][1] ), .B(
        \u_div/SumTmp[49][1] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_50_1  ( .A(\u_div/SumTmp[50][1] ), .B(
        \u_div/SumTmp[50][1] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_52_1  ( .A(\u_div/SumTmp[52][1] ), .B(
        \u_div/SumTmp[52][1] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_53_1  ( .A(\u_div/SumTmp[53][1] ), .B(
        \u_div/SumTmp[53][1] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_1_3  ( .A(\u_div/PartRem[2][3] ), .B(
        \u_div/SumTmp[1][3] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_3  ( .A(\u_div/PartRem[3][3] ), .B(
        \u_div/SumTmp[2][3] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_1_4  ( .A(\u_div/PartRem[2][4] ), .B(
        \u_div/SumTmp[1][4] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_4  ( .A(\u_div/PartRem[4][4] ), .B(
        \u_div/SumTmp[3][4] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_4  ( .A(\u_div/PartRem[3][4] ), .B(
        \u_div/SumTmp[2][4] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_4  ( .A(\u_div/PartRem[5][4] ), .B(
        \u_div/SumTmp[4][4] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_4  ( .A(\u_div/PartRem[6][4] ), .B(
        \u_div/SumTmp[5][4] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_9_4  ( .A(\u_div/PartRem[10][4] ), .B(
        \u_div/SumTmp[9][4] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_4  ( .A(\u_div/PartRem[7][4] ), .B(
        \u_div/SumTmp[6][4] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_4  ( .A(\u_div/PartRem[11][4] ), .B(
        \u_div/SumTmp[10][4] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_8_4  ( .A(\u_div/PartRem[9][4] ), .B(
        \u_div/SumTmp[8][4] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_4  ( .A(\u_div/PartRem[8][4] ), .B(
        \u_div/SumTmp[7][4] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_4  ( .A(\u_div/PartRem[23][4] ), .B(
        \u_div/SumTmp[22][4] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_4  ( .A(\u_div/PartRem[12][4] ), .B(
        \u_div/SumTmp[11][4] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_4  ( .A(\u_div/PartRem[21][4] ), .B(
        \u_div/SumTmp[20][4] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_4  ( .A(\u_div/PartRem[26][4] ), .B(
        \u_div/SumTmp[25][4] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_4  ( .A(\u_div/PartRem[13][4] ), .B(
        \u_div/SumTmp[12][4] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_4  ( .A(\u_div/PartRem[22][4] ), .B(
        \u_div/SumTmp[21][4] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_4  ( .A(\u_div/PartRem[25][4] ), .B(
        \u_div/SumTmp[24][4] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_4  ( .A(\u_div/PartRem[24][4] ), .B(
        \u_div/SumTmp[23][4] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_4  ( .A(\u_div/PartRem[14][4] ), .B(
        \u_div/SumTmp[13][4] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_4  ( .A(\u_div/PartRem[20][4] ), .B(
        \u_div/SumTmp[19][4] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_4  ( .A(\u_div/PartRem[15][4] ), .B(
        \u_div/SumTmp[14][4] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_4  ( .A(\u_div/PartRem[29][4] ), .B(
        \u_div/SumTmp[28][4] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_4  ( .A(\u_div/PartRem[16][4] ), .B(
        \u_div/SumTmp[15][4] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_4  ( .A(\u_div/PartRem[19][4] ), .B(
        \u_div/SumTmp[18][4] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_4  ( .A(\u_div/PartRem[17][4] ), .B(
        \u_div/SumTmp[16][4] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_4  ( .A(\u_div/PartRem[18][4] ), .B(
        \u_div/SumTmp[17][4] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_4  ( .A(\u_div/PartRem[27][4] ), .B(
        \u_div/SumTmp[26][4] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_4  ( .A(\u_div/PartRem[28][4] ), .B(
        \u_div/SumTmp[27][4] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_4  ( .A(\u_div/PartRem[30][4] ), .B(
        \u_div/SumTmp[29][4] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_4  ( .A(\u_div/PartRem[31][4] ), .B(
        \u_div/SumTmp[30][4] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_4  ( .A(\u_div/PartRem[34][4] ), .B(
        \u_div/SumTmp[33][4] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_4  ( .A(\u_div/PartRem[32][4] ), .B(
        \u_div/SumTmp[31][4] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_4  ( .A(\u_div/PartRem[33][4] ), .B(
        \u_div/SumTmp[32][4] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_4  ( .A(\u_div/PartRem[35][4] ), .B(
        \u_div/SumTmp[34][4] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_4  ( .A(\u_div/PartRem[36][4] ), .B(
        \u_div/SumTmp[35][4] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_4  ( .A(\u_div/PartRem[39][4] ), .B(
        \u_div/SumTmp[38][4] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_4  ( .A(\u_div/PartRem[37][4] ), .B(
        \u_div/SumTmp[36][4] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_4  ( .A(\u_div/PartRem[38][4] ), .B(
        \u_div/SumTmp[37][4] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_4  ( .A(\u_div/PartRem[40][4] ), .B(
        \u_div/SumTmp[39][4] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_4  ( .A(\u_div/PartRem[41][4] ), .B(
        \u_div/SumTmp[40][4] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_4  ( .A(\u_div/PartRem[44][4] ), .B(
        \u_div/SumTmp[43][4] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_4  ( .A(\u_div/PartRem[42][4] ), .B(
        \u_div/SumTmp[41][4] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_4  ( .A(\u_div/PartRem[47][4] ), .B(
        \u_div/SumTmp[46][4] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_4  ( .A(\u_div/PartRem[43][4] ), .B(
        \u_div/SumTmp[42][4] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_4  ( .A(\u_div/PartRem[50][4] ), .B(
        \u_div/SumTmp[49][4] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_4  ( .A(\u_div/PartRem[52][4] ), .B(
        \u_div/SumTmp[51][4] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_4  ( .A(\u_div/PartRem[46][4] ), .B(
        \u_div/SumTmp[45][4] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_4  ( .A(\u_div/PartRem[45][4] ), .B(
        \u_div/SumTmp[44][4] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_4  ( .A(\u_div/PartRem[49][4] ), .B(
        \u_div/SumTmp[48][4] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_4  ( .A(\u_div/PartRem[55][4] ), .B(
        \u_div/SumTmp[54][4] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_4  ( .A(\u_div/PartRem[51][4] ), .B(
        \u_div/SumTmp[50][4] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_4  ( .A(\u_div/PartRem[48][4] ), .B(
        \u_div/SumTmp[47][4] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_4  ( .A(\u_div/PartRem[54][4] ), .B(
        \u_div/SumTmp[53][4] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_4  ( .A(\u_div/PartRem[53][4] ), .B(
        \u_div/SumTmp[52][4] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_4  ( .A(\u_div/PartRem[58][4] ), .B(
        \u_div/SumTmp[57][4] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_4  ( .A(\u_div/PartRem[56][4] ), .B(
        \u_div/SumTmp[55][4] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_4  ( .A(\u_div/PartRem[57][4] ), .B(
        \u_div/SumTmp[56][4] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_4  ( .A(\u_div/PartRem[59][4] ), .B(
        \u_div/SumTmp[58][4] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][5] ) );
  MX2X2 \u_div/u_mx_PartRem_1_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/SumTmp[1][2] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][3] ) );
  CLKMX2X8 \u_div/u_mx_PartRem_1_3_1  ( .A(\u_div/SumTmp[3][1] ), .B(
        \u_div/SumTmp[3][1] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][2] ) );
  ADDHX1 U1 ( .A(\u_div/PartRem[8][4] ), .B(\u_div/u_add_PartRem_2_7/n3 ), 
        .CO(\u_div/u_add_PartRem_2_7/n2 ), .S(\u_div/SumTmp[7][4] ) );
  XOR2XL U2 ( .A(\u_div/CryTmp[3][6] ), .B(n3), .Y(\u_div/QInv[3] ) );
  MXI2X2 U3 ( .A(\u_div/SumTmp[3][2] ), .B(\u_div/PartRem[4][2] ), .S0(
        \u_div/CryTmp[3][6] ), .Y(\u_div/PartRem[3][3] ) );
  OR2X6 U4 ( .A(\u_div/PartRem[4][5] ), .B(\u_div/u_add_PartRem_2_3/n2 ), .Y(
        \u_div/CryTmp[3][6] ) );
  INVX3 U5 ( .A(\u_div/QInv[63] ), .Y(n2) );
  OR2X1 U6 ( .A(\u_div/PartRem[13][2] ), .B(\u_div/PartRem[13][3] ), .Y(
        \u_div/u_add_PartRem_2_12/n3 ) );
  OR2X1 U7 ( .A(\u_div/PartRem[18][2] ), .B(\u_div/PartRem[18][3] ), .Y(
        \u_div/u_add_PartRem_2_17/n3 ) );
  OR2X1 U8 ( .A(\u_div/PartRem[23][2] ), .B(\u_div/PartRem[23][3] ), .Y(
        \u_div/u_add_PartRem_2_22/n3 ) );
  OR2X1 U9 ( .A(\u_div/PartRem[8][2] ), .B(\u_div/PartRem[8][3] ), .Y(
        \u_div/u_add_PartRem_2_7/n3 ) );
  OR2X1 U10 ( .A(\u_div/PartRem[28][2] ), .B(\u_div/PartRem[28][3] ), .Y(
        \u_div/u_add_PartRem_2_27/n3 ) );
  OR2X1 U11 ( .A(\u_div/PartRem[33][2] ), .B(\u_div/PartRem[33][3] ), .Y(
        \u_div/u_add_PartRem_2_32/n3 ) );
  OR2X1 U12 ( .A(\u_div/PartRem[38][2] ), .B(\u_div/PartRem[38][3] ), .Y(
        \u_div/u_add_PartRem_2_37/n3 ) );
  OR2X1 U13 ( .A(\u_div/PartRem[43][2] ), .B(\u_div/PartRem[43][3] ), .Y(
        \u_div/u_add_PartRem_2_42/n3 ) );
  OR2X1 U14 ( .A(\u_div/PartRem[48][2] ), .B(\u_div/PartRem[48][3] ), .Y(
        \u_div/u_add_PartRem_2_47/n3 ) );
  OR2X1 U15 ( .A(\u_div/PartRem[53][2] ), .B(\u_div/PartRem[53][3] ), .Y(
        \u_div/u_add_PartRem_2_52/n3 ) );
  OR2X2 U16 ( .A(\u_div/PartRem[54][2] ), .B(\u_div/PartRem[54][3] ), .Y(
        \u_div/u_add_PartRem_2_53/n3 ) );
  OR2X2 U17 ( .A(\u_div/PartRem[55][2] ), .B(\u_div/PartRem[55][3] ), .Y(
        \u_div/u_add_PartRem_2_54/n3 ) );
  OR2X2 U18 ( .A(\u_div/PartRem[56][2] ), .B(\u_div/PartRem[56][3] ), .Y(
        \u_div/u_add_PartRem_2_55/n3 ) );
  OR2X2 U19 ( .A(\u_div/PartRem[57][2] ), .B(\u_div/PartRem[57][3] ), .Y(
        \u_div/u_add_PartRem_2_56/n3 ) );
  OR2X2 U20 ( .A(\u_div/PartRem[58][2] ), .B(\u_div/PartRem[58][3] ), .Y(
        \u_div/u_add_PartRem_2_57/n3 ) );
  NOR2X2 U21 ( .A(\u_div/PartRem[63][0] ), .B(\u_div/PartRem[62][0] ), .Y(n8)
         );
  OR2X6 U22 ( .A(\u_div/PartRem[3][5] ), .B(\u_div/u_add_PartRem_2_2/n2 ), .Y(
        \u_div/CryTmp[2][6] ) );
  NOR2BX4 U23 ( .AN(\u_div/PartRem[64][0] ), .B(n8), .Y(\u_div/CryTmp[59][6] )
         );
  XOR2X4 U24 ( .A(\u_div/CryTmp[0][6] ), .B(n5), .Y(\u_div/QInv[0] ) );
  AO21X4 U25 ( .A0(\u_div/PartRem[1][4] ), .A1(n6), .B0(\u_div/PartRem[1][5] ), 
        .Y(\u_div/CryTmp[0][6] ) );
  OR2X1 U26 ( .A(\u_div/PartRem[4][2] ), .B(\u_div/PartRem[4][3] ), .Y(
        \u_div/u_add_PartRem_2_3/n3 ) );
  ADDHX1 U27 ( .A(\u_div/PartRem[2][4] ), .B(\u_div/u_add_PartRem_2_1/n3 ), 
        .CO(\u_div/u_add_PartRem_2_1/n2 ), .S(\u_div/SumTmp[1][4] ) );
  XNOR2XL U28 ( .A(\u_div/PartRem[64][0] ), .B(n8), .Y(\u_div/SumTmp[59][4] )
         );
  OR2X6 U29 ( .A(\u_div/PartRem[2][5] ), .B(\u_div/u_add_PartRem_2_1/n2 ), .Y(
        \u_div/CryTmp[1][6] ) );
  XOR2XL U30 ( .A(\u_div/CryTmp[51][6] ), .B(n4), .Y(\u_div/QInv[51] ) );
  XOR2XL U31 ( .A(\u_div/CryTmp[52][6] ), .B(n5), .Y(\u_div/QInv[52] ) );
  XOR2XL U32 ( .A(\u_div/CryTmp[41][6] ), .B(n5), .Y(\u_div/QInv[41] ) );
  XOR2XL U33 ( .A(\u_div/CryTmp[31][6] ), .B(n5), .Y(\u_div/QInv[31] ) );
  XOR2XL U34 ( .A(\u_div/CryTmp[11][6] ), .B(n4), .Y(\u_div/QInv[11] ) );
  XOR2XL U35 ( .A(\u_div/CryTmp[12][6] ), .B(n5), .Y(\u_div/QInv[12] ) );
  XOR2XL U36 ( .A(\u_div/CryTmp[1][6] ), .B(n4), .Y(\u_div/QInv[1] ) );
  XOR2XL U37 ( .A(\u_div/CryTmp[22][6] ), .B(n4), .Y(\u_div/QInv[22] ) );
  XOR2XL U38 ( .A(\u_div/CryTmp[32][6] ), .B(n3), .Y(\u_div/QInv[32] ) );
  XOR2XL U39 ( .A(\u_div/CryTmp[21][6] ), .B(n3), .Y(\u_div/QInv[21] ) );
  INVXL U40 ( .A(\u_div/PartRem[59][2] ), .Y(\u_div/SumTmp[58][2] ) );
  INVXL U41 ( .A(\u_div/PartRem[58][2] ), .Y(\u_div/SumTmp[57][2] ) );
  INVXL U42 ( .A(\u_div/PartRem[57][2] ), .Y(\u_div/SumTmp[56][2] ) );
  INVXL U43 ( .A(\u_div/PartRem[56][2] ), .Y(\u_div/SumTmp[55][2] ) );
  INVXL U44 ( .A(\u_div/PartRem[55][2] ), .Y(\u_div/SumTmp[54][2] ) );
  INVXL U45 ( .A(\u_div/PartRem[54][2] ), .Y(\u_div/SumTmp[53][2] ) );
  INVX3 U46 ( .A(n2), .Y(n3) );
  ADDHX2 U47 ( .A(\u_div/PartRem[3][4] ), .B(\u_div/u_add_PartRem_2_2/n3 ), 
        .CO(\u_div/u_add_PartRem_2_2/n2 ), .S(\u_div/SumTmp[2][4] ) );
  OR2X2 U48 ( .A(\u_div/PartRem[3][2] ), .B(\u_div/PartRem[3][3] ), .Y(
        \u_div/u_add_PartRem_2_2/n3 ) );
  ADDHX2 U49 ( .A(\u_div/PartRem[59][4] ), .B(\u_div/u_add_PartRem_2_58/n3 ), 
        .CO(\u_div/u_add_PartRem_2_58/n2 ), .S(\u_div/SumTmp[58][4] ) );
  OR2X6 U50 ( .A(\u_div/PartRem[59][2] ), .B(\u_div/PartRem[59][3] ), .Y(
        \u_div/u_add_PartRem_2_58/n3 ) );
  ADDHX2 U51 ( .A(\u_div/PartRem[55][4] ), .B(\u_div/u_add_PartRem_2_54/n3 ), 
        .CO(\u_div/u_add_PartRem_2_54/n2 ), .S(\u_div/SumTmp[54][4] ) );
  ADDHX2 U52 ( .A(\u_div/PartRem[54][4] ), .B(\u_div/u_add_PartRem_2_53/n3 ), 
        .CO(\u_div/u_add_PartRem_2_53/n2 ), .S(\u_div/SumTmp[53][4] ) );
  ADDHX2 U53 ( .A(\u_div/PartRem[52][4] ), .B(\u_div/u_add_PartRem_2_51/n3 ), 
        .CO(\u_div/u_add_PartRem_2_51/n2 ), .S(\u_div/SumTmp[51][4] ) );
  OR2X2 U54 ( .A(\u_div/PartRem[52][2] ), .B(\u_div/PartRem[52][3] ), .Y(
        \u_div/u_add_PartRem_2_51/n3 ) );
  ADDHX2 U55 ( .A(\u_div/PartRem[45][4] ), .B(\u_div/u_add_PartRem_2_44/n3 ), 
        .CO(\u_div/u_add_PartRem_2_44/n2 ), .S(\u_div/SumTmp[44][4] ) );
  OR2X2 U56 ( .A(\u_div/PartRem[45][2] ), .B(\u_div/PartRem[45][3] ), .Y(
        \u_div/u_add_PartRem_2_44/n3 ) );
  ADDHX2 U57 ( .A(\u_div/PartRem[51][4] ), .B(\u_div/u_add_PartRem_2_50/n3 ), 
        .CO(\u_div/u_add_PartRem_2_50/n2 ), .S(\u_div/SumTmp[50][4] ) );
  OR2X2 U58 ( .A(\u_div/PartRem[51][2] ), .B(\u_div/PartRem[51][3] ), .Y(
        \u_div/u_add_PartRem_2_50/n3 ) );
  ADDHX2 U59 ( .A(\u_div/PartRem[50][4] ), .B(\u_div/u_add_PartRem_2_49/n3 ), 
        .CO(\u_div/u_add_PartRem_2_49/n2 ), .S(\u_div/SumTmp[49][4] ) );
  OR2X2 U60 ( .A(\u_div/PartRem[50][2] ), .B(\u_div/PartRem[50][3] ), .Y(
        \u_div/u_add_PartRem_2_49/n3 ) );
  ADDHX2 U61 ( .A(\u_div/PartRem[49][4] ), .B(\u_div/u_add_PartRem_2_48/n3 ), 
        .CO(\u_div/u_add_PartRem_2_48/n2 ), .S(\u_div/SumTmp[48][4] ) );
  OR2X2 U62 ( .A(\u_div/PartRem[49][2] ), .B(\u_div/PartRem[49][3] ), .Y(
        \u_div/u_add_PartRem_2_48/n3 ) );
  ADDHX2 U63 ( .A(\u_div/PartRem[47][4] ), .B(\u_div/u_add_PartRem_2_46/n3 ), 
        .CO(\u_div/u_add_PartRem_2_46/n2 ), .S(\u_div/SumTmp[46][4] ) );
  OR2X2 U64 ( .A(\u_div/PartRem[47][2] ), .B(\u_div/PartRem[47][3] ), .Y(
        \u_div/u_add_PartRem_2_46/n3 ) );
  ADDHX2 U65 ( .A(\u_div/PartRem[46][4] ), .B(\u_div/u_add_PartRem_2_45/n3 ), 
        .CO(\u_div/u_add_PartRem_2_45/n2 ), .S(\u_div/SumTmp[45][4] ) );
  OR2X2 U66 ( .A(\u_div/PartRem[46][2] ), .B(\u_div/PartRem[46][3] ), .Y(
        \u_div/u_add_PartRem_2_45/n3 ) );
  ADDHX2 U67 ( .A(\u_div/PartRem[44][4] ), .B(\u_div/u_add_PartRem_2_43/n3 ), 
        .CO(\u_div/u_add_PartRem_2_43/n2 ), .S(\u_div/SumTmp[43][4] ) );
  OR2X2 U68 ( .A(\u_div/PartRem[44][2] ), .B(\u_div/PartRem[44][3] ), .Y(
        \u_div/u_add_PartRem_2_43/n3 ) );
  ADDHX2 U69 ( .A(\u_div/PartRem[42][4] ), .B(\u_div/u_add_PartRem_2_41/n3 ), 
        .CO(\u_div/u_add_PartRem_2_41/n2 ), .S(\u_div/SumTmp[41][4] ) );
  OR2X2 U70 ( .A(\u_div/PartRem[42][2] ), .B(\u_div/PartRem[42][3] ), .Y(
        \u_div/u_add_PartRem_2_41/n3 ) );
  ADDHX2 U71 ( .A(\u_div/PartRem[41][4] ), .B(\u_div/u_add_PartRem_2_40/n3 ), 
        .CO(\u_div/u_add_PartRem_2_40/n2 ), .S(\u_div/SumTmp[40][4] ) );
  OR2X2 U72 ( .A(\u_div/PartRem[41][2] ), .B(\u_div/PartRem[41][3] ), .Y(
        \u_div/u_add_PartRem_2_40/n3 ) );
  ADDHX2 U73 ( .A(\u_div/PartRem[40][4] ), .B(\u_div/u_add_PartRem_2_39/n3 ), 
        .CO(\u_div/u_add_PartRem_2_39/n2 ), .S(\u_div/SumTmp[39][4] ) );
  OR2X2 U74 ( .A(\u_div/PartRem[40][2] ), .B(\u_div/PartRem[40][3] ), .Y(
        \u_div/u_add_PartRem_2_39/n3 ) );
  ADDHX2 U75 ( .A(\u_div/PartRem[39][4] ), .B(\u_div/u_add_PartRem_2_38/n3 ), 
        .CO(\u_div/u_add_PartRem_2_38/n2 ), .S(\u_div/SumTmp[38][4] ) );
  OR2X2 U76 ( .A(\u_div/PartRem[39][2] ), .B(\u_div/PartRem[39][3] ), .Y(
        \u_div/u_add_PartRem_2_38/n3 ) );
  ADDHX2 U77 ( .A(\u_div/PartRem[37][4] ), .B(\u_div/u_add_PartRem_2_36/n3 ), 
        .CO(\u_div/u_add_PartRem_2_36/n2 ), .S(\u_div/SumTmp[36][4] ) );
  OR2X2 U78 ( .A(\u_div/PartRem[37][2] ), .B(\u_div/PartRem[37][3] ), .Y(
        \u_div/u_add_PartRem_2_36/n3 ) );
  ADDHX2 U79 ( .A(\u_div/PartRem[36][4] ), .B(\u_div/u_add_PartRem_2_35/n3 ), 
        .CO(\u_div/u_add_PartRem_2_35/n2 ), .S(\u_div/SumTmp[35][4] ) );
  OR2X2 U80 ( .A(\u_div/PartRem[36][2] ), .B(\u_div/PartRem[36][3] ), .Y(
        \u_div/u_add_PartRem_2_35/n3 ) );
  ADDHX2 U81 ( .A(\u_div/PartRem[35][4] ), .B(\u_div/u_add_PartRem_2_34/n3 ), 
        .CO(\u_div/u_add_PartRem_2_34/n2 ), .S(\u_div/SumTmp[34][4] ) );
  OR2X2 U82 ( .A(\u_div/PartRem[35][2] ), .B(\u_div/PartRem[35][3] ), .Y(
        \u_div/u_add_PartRem_2_34/n3 ) );
  ADDHX2 U83 ( .A(\u_div/PartRem[34][4] ), .B(\u_div/u_add_PartRem_2_33/n3 ), 
        .CO(\u_div/u_add_PartRem_2_33/n2 ), .S(\u_div/SumTmp[33][4] ) );
  OR2X2 U84 ( .A(\u_div/PartRem[34][2] ), .B(\u_div/PartRem[34][3] ), .Y(
        \u_div/u_add_PartRem_2_33/n3 ) );
  ADDHX2 U85 ( .A(\u_div/PartRem[32][4] ), .B(\u_div/u_add_PartRem_2_31/n3 ), 
        .CO(\u_div/u_add_PartRem_2_31/n2 ), .S(\u_div/SumTmp[31][4] ) );
  OR2X2 U86 ( .A(\u_div/PartRem[32][2] ), .B(\u_div/PartRem[32][3] ), .Y(
        \u_div/u_add_PartRem_2_31/n3 ) );
  ADDHX2 U87 ( .A(\u_div/PartRem[31][4] ), .B(\u_div/u_add_PartRem_2_30/n3 ), 
        .CO(\u_div/u_add_PartRem_2_30/n2 ), .S(\u_div/SumTmp[30][4] ) );
  OR2X2 U88 ( .A(\u_div/PartRem[31][2] ), .B(\u_div/PartRem[31][3] ), .Y(
        \u_div/u_add_PartRem_2_30/n3 ) );
  ADDHX2 U89 ( .A(\u_div/PartRem[30][4] ), .B(\u_div/u_add_PartRem_2_29/n3 ), 
        .CO(\u_div/u_add_PartRem_2_29/n2 ), .S(\u_div/SumTmp[29][4] ) );
  OR2X2 U90 ( .A(\u_div/PartRem[30][2] ), .B(\u_div/PartRem[30][3] ), .Y(
        \u_div/u_add_PartRem_2_29/n3 ) );
  ADDHX2 U91 ( .A(\u_div/PartRem[29][4] ), .B(\u_div/u_add_PartRem_2_28/n3 ), 
        .CO(\u_div/u_add_PartRem_2_28/n2 ), .S(\u_div/SumTmp[28][4] ) );
  OR2X2 U92 ( .A(\u_div/PartRem[29][2] ), .B(\u_div/PartRem[29][3] ), .Y(
        \u_div/u_add_PartRem_2_28/n3 ) );
  ADDHX2 U93 ( .A(\u_div/PartRem[27][4] ), .B(\u_div/u_add_PartRem_2_26/n3 ), 
        .CO(\u_div/u_add_PartRem_2_26/n2 ), .S(\u_div/SumTmp[26][4] ) );
  OR2X2 U94 ( .A(\u_div/PartRem[27][2] ), .B(\u_div/PartRem[27][3] ), .Y(
        \u_div/u_add_PartRem_2_26/n3 ) );
  ADDHX2 U95 ( .A(\u_div/PartRem[17][4] ), .B(\u_div/u_add_PartRem_2_16/n3 ), 
        .CO(\u_div/u_add_PartRem_2_16/n2 ), .S(\u_div/SumTmp[16][4] ) );
  OR2X2 U96 ( .A(\u_div/PartRem[17][2] ), .B(\u_div/PartRem[17][3] ), .Y(
        \u_div/u_add_PartRem_2_16/n3 ) );
  ADDHX2 U97 ( .A(\u_div/PartRem[16][4] ), .B(\u_div/u_add_PartRem_2_15/n3 ), 
        .CO(\u_div/u_add_PartRem_2_15/n2 ), .S(\u_div/SumTmp[15][4] ) );
  OR2X2 U98 ( .A(\u_div/PartRem[16][2] ), .B(\u_div/PartRem[16][3] ), .Y(
        \u_div/u_add_PartRem_2_15/n3 ) );
  ADDHX2 U99 ( .A(\u_div/PartRem[15][4] ), .B(\u_div/u_add_PartRem_2_14/n3 ), 
        .CO(\u_div/u_add_PartRem_2_14/n2 ), .S(\u_div/SumTmp[14][4] ) );
  OR2X2 U100 ( .A(\u_div/PartRem[15][2] ), .B(\u_div/PartRem[15][3] ), .Y(
        \u_div/u_add_PartRem_2_14/n3 ) );
  ADDHX2 U101 ( .A(\u_div/PartRem[19][4] ), .B(\u_div/u_add_PartRem_2_18/n3 ), 
        .CO(\u_div/u_add_PartRem_2_18/n2 ), .S(\u_div/SumTmp[18][4] ) );
  OR2X2 U102 ( .A(\u_div/PartRem[19][2] ), .B(\u_div/PartRem[19][3] ), .Y(
        \u_div/u_add_PartRem_2_18/n3 ) );
  ADDHX2 U103 ( .A(\u_div/PartRem[14][4] ), .B(\u_div/u_add_PartRem_2_13/n3 ), 
        .CO(\u_div/u_add_PartRem_2_13/n2 ), .S(\u_div/SumTmp[13][4] ) );
  OR2X2 U104 ( .A(\u_div/PartRem[14][2] ), .B(\u_div/PartRem[14][3] ), .Y(
        \u_div/u_add_PartRem_2_13/n3 ) );
  ADDHX2 U105 ( .A(\u_div/PartRem[26][4] ), .B(\u_div/u_add_PartRem_2_25/n3 ), 
        .CO(\u_div/u_add_PartRem_2_25/n2 ), .S(\u_div/SumTmp[25][4] ) );
  OR2X2 U106 ( .A(\u_div/PartRem[26][2] ), .B(\u_div/PartRem[26][3] ), .Y(
        \u_div/u_add_PartRem_2_25/n3 ) );
  ADDHX2 U107 ( .A(\u_div/PartRem[24][4] ), .B(\u_div/u_add_PartRem_2_23/n3 ), 
        .CO(\u_div/u_add_PartRem_2_23/n2 ), .S(\u_div/SumTmp[23][4] ) );
  OR2X2 U108 ( .A(\u_div/PartRem[24][2] ), .B(\u_div/PartRem[24][3] ), .Y(
        \u_div/u_add_PartRem_2_23/n3 ) );
  ADDHX2 U109 ( .A(\u_div/PartRem[25][4] ), .B(\u_div/u_add_PartRem_2_24/n3 ), 
        .CO(\u_div/u_add_PartRem_2_24/n2 ), .S(\u_div/SumTmp[24][4] ) );
  OR2X2 U110 ( .A(\u_div/PartRem[25][2] ), .B(\u_div/PartRem[25][3] ), .Y(
        \u_div/u_add_PartRem_2_24/n3 ) );
  ADDHX2 U111 ( .A(\u_div/PartRem[20][4] ), .B(\u_div/u_add_PartRem_2_19/n3 ), 
        .CO(\u_div/u_add_PartRem_2_19/n2 ), .S(\u_div/SumTmp[19][4] ) );
  OR2X2 U112 ( .A(\u_div/PartRem[20][2] ), .B(\u_div/PartRem[20][3] ), .Y(
        \u_div/u_add_PartRem_2_19/n3 ) );
  ADDHX2 U113 ( .A(\u_div/PartRem[21][4] ), .B(\u_div/u_add_PartRem_2_20/n3 ), 
        .CO(\u_div/u_add_PartRem_2_20/n2 ), .S(\u_div/SumTmp[20][4] ) );
  OR2X2 U114 ( .A(\u_div/PartRem[21][2] ), .B(\u_div/PartRem[21][3] ), .Y(
        \u_div/u_add_PartRem_2_20/n3 ) );
  ADDHX2 U115 ( .A(\u_div/PartRem[12][4] ), .B(\u_div/u_add_PartRem_2_11/n3 ), 
        .CO(\u_div/u_add_PartRem_2_11/n2 ), .S(\u_div/SumTmp[11][4] ) );
  OR2X2 U116 ( .A(\u_div/PartRem[12][2] ), .B(\u_div/PartRem[12][3] ), .Y(
        \u_div/u_add_PartRem_2_11/n3 ) );
  ADDHX2 U117 ( .A(\u_div/PartRem[22][4] ), .B(\u_div/u_add_PartRem_2_21/n3 ), 
        .CO(\u_div/u_add_PartRem_2_21/n2 ), .S(\u_div/SumTmp[21][4] ) );
  OR2X2 U118 ( .A(\u_div/PartRem[22][2] ), .B(\u_div/PartRem[22][3] ), .Y(
        \u_div/u_add_PartRem_2_21/n3 ) );
  ADDHX2 U119 ( .A(\u_div/PartRem[11][4] ), .B(\u_div/u_add_PartRem_2_10/n3 ), 
        .CO(\u_div/u_add_PartRem_2_10/n2 ), .S(\u_div/SumTmp[10][4] ) );
  OR2X2 U120 ( .A(\u_div/PartRem[11][2] ), .B(\u_div/PartRem[11][3] ), .Y(
        \u_div/u_add_PartRem_2_10/n3 ) );
  ADDHX2 U121 ( .A(\u_div/PartRem[7][4] ), .B(\u_div/u_add_PartRem_2_6/n3 ), 
        .CO(\u_div/u_add_PartRem_2_6/n2 ), .S(\u_div/SumTmp[6][4] ) );
  OR2X2 U122 ( .A(\u_div/PartRem[7][2] ), .B(\u_div/PartRem[7][3] ), .Y(
        \u_div/u_add_PartRem_2_6/n3 ) );
  ADDHX2 U123 ( .A(\u_div/PartRem[9][4] ), .B(\u_div/u_add_PartRem_2_8/n3 ), 
        .CO(\u_div/u_add_PartRem_2_8/n2 ), .S(\u_div/SumTmp[8][4] ) );
  OR2X2 U124 ( .A(\u_div/PartRem[9][2] ), .B(\u_div/PartRem[9][3] ), .Y(
        \u_div/u_add_PartRem_2_8/n3 ) );
  ADDHX2 U125 ( .A(\u_div/PartRem[10][4] ), .B(\u_div/u_add_PartRem_2_9/n3 ), 
        .CO(\u_div/u_add_PartRem_2_9/n2 ), .S(\u_div/SumTmp[9][4] ) );
  OR2X2 U126 ( .A(\u_div/PartRem[10][2] ), .B(\u_div/PartRem[10][3] ), .Y(
        \u_div/u_add_PartRem_2_9/n3 ) );
  ADDHX2 U127 ( .A(\u_div/PartRem[6][4] ), .B(\u_div/u_add_PartRem_2_5/n3 ), 
        .CO(\u_div/u_add_PartRem_2_5/n2 ), .S(\u_div/SumTmp[5][4] ) );
  OR2X2 U128 ( .A(\u_div/PartRem[6][2] ), .B(\u_div/PartRem[6][3] ), .Y(
        \u_div/u_add_PartRem_2_5/n3 ) );
  ADDHX2 U129 ( .A(\u_div/PartRem[5][4] ), .B(\u_div/u_add_PartRem_2_4/n3 ), 
        .CO(\u_div/u_add_PartRem_2_4/n2 ), .S(\u_div/SumTmp[4][4] ) );
  OR2X2 U130 ( .A(\u_div/PartRem[5][2] ), .B(\u_div/PartRem[5][3] ), .Y(
        \u_div/u_add_PartRem_2_4/n3 ) );
  OR2X2 U131 ( .A(\u_div/PartRem[2][2] ), .B(\u_div/PartRem[2][3] ), .Y(
        \u_div/u_add_PartRem_2_1/n3 ) );
  ADDHX2 U132 ( .A(\u_div/PartRem[58][4] ), .B(\u_div/u_add_PartRem_2_57/n3 ), 
        .CO(\u_div/u_add_PartRem_2_57/n2 ), .S(\u_div/SumTmp[57][4] ) );
  ADDHX2 U133 ( .A(\u_div/PartRem[56][4] ), .B(\u_div/u_add_PartRem_2_55/n3 ), 
        .CO(\u_div/u_add_PartRem_2_55/n2 ), .S(\u_div/SumTmp[55][4] ) );
  ADDHX2 U134 ( .A(\u_div/PartRem[57][4] ), .B(\u_div/u_add_PartRem_2_56/n3 ), 
        .CO(\u_div/u_add_PartRem_2_56/n2 ), .S(\u_div/SumTmp[56][4] ) );
  MXI2X1 U135 ( .A(\u_div/SumTmp[1][1] ), .B(\u_div/SumTmp[1][1] ), .S0(
        \u_div/CryTmp[1][6] ), .Y(n1) );
  INVXL U136 ( .A(\u_div/PartRem[2][2] ), .Y(\u_div/SumTmp[1][2] ) );
  CLKINVX1 U137 ( .A(\u_div/PartRem[4][2] ), .Y(\u_div/SumTmp[3][2] ) );
  MXI2X1 U138 ( .A(n7), .B(\u_div/PartRem[62][0] ), .S0(\u_div/CryTmp[59][6] ), 
        .Y(\u_div/PartRem[59][3] ) );
  CLKINVX1 U139 ( .A(\u_div/PartRem[62][0] ), .Y(n7) );
  MXI2X1 U140 ( .A(\u_div/SumTmp[4][2] ), .B(\u_div/PartRem[5][2] ), .S0(
        \u_div/CryTmp[4][6] ), .Y(\u_div/PartRem[4][3] ) );
  CLKINVX1 U141 ( .A(\u_div/PartRem[5][2] ), .Y(\u_div/SumTmp[4][2] ) );
  MXI2X1 U142 ( .A(\u_div/SumTmp[53][2] ), .B(\u_div/PartRem[54][2] ), .S0(
        \u_div/CryTmp[53][6] ), .Y(\u_div/PartRem[53][3] ) );
  MXI2X1 U143 ( .A(\u_div/SumTmp[48][2] ), .B(\u_div/PartRem[49][2] ), .S0(
        \u_div/CryTmp[48][6] ), .Y(\u_div/PartRem[48][3] ) );
  CLKINVX1 U144 ( .A(\u_div/PartRem[49][2] ), .Y(\u_div/SumTmp[48][2] ) );
  MXI2X1 U145 ( .A(\u_div/SumTmp[43][2] ), .B(\u_div/PartRem[44][2] ), .S0(
        \u_div/CryTmp[43][6] ), .Y(\u_div/PartRem[43][3] ) );
  CLKINVX1 U146 ( .A(\u_div/PartRem[44][2] ), .Y(\u_div/SumTmp[43][2] ) );
  MXI2X1 U147 ( .A(\u_div/SumTmp[38][2] ), .B(\u_div/PartRem[39][2] ), .S0(
        \u_div/CryTmp[38][6] ), .Y(\u_div/PartRem[38][3] ) );
  CLKINVX1 U148 ( .A(\u_div/PartRem[39][2] ), .Y(\u_div/SumTmp[38][2] ) );
  MXI2X1 U149 ( .A(\u_div/SumTmp[33][2] ), .B(\u_div/PartRem[34][2] ), .S0(
        \u_div/CryTmp[33][6] ), .Y(\u_div/PartRem[33][3] ) );
  CLKINVX1 U150 ( .A(\u_div/PartRem[34][2] ), .Y(\u_div/SumTmp[33][2] ) );
  MXI2X1 U151 ( .A(\u_div/SumTmp[28][2] ), .B(\u_div/PartRem[29][2] ), .S0(
        \u_div/CryTmp[28][6] ), .Y(\u_div/PartRem[28][3] ) );
  CLKINVX1 U152 ( .A(\u_div/PartRem[29][2] ), .Y(\u_div/SumTmp[28][2] ) );
  MXI2X1 U153 ( .A(\u_div/SumTmp[23][2] ), .B(\u_div/PartRem[24][2] ), .S0(
        \u_div/CryTmp[23][6] ), .Y(\u_div/PartRem[23][3] ) );
  CLKINVX1 U154 ( .A(\u_div/PartRem[24][2] ), .Y(\u_div/SumTmp[23][2] ) );
  MXI2X1 U155 ( .A(\u_div/SumTmp[18][2] ), .B(\u_div/PartRem[19][2] ), .S0(
        \u_div/CryTmp[18][6] ), .Y(\u_div/PartRem[18][3] ) );
  CLKINVX1 U156 ( .A(\u_div/PartRem[19][2] ), .Y(\u_div/SumTmp[18][2] ) );
  MXI2X1 U157 ( .A(\u_div/SumTmp[13][2] ), .B(\u_div/PartRem[14][2] ), .S0(
        \u_div/CryTmp[13][6] ), .Y(\u_div/PartRem[13][3] ) );
  CLKINVX1 U158 ( .A(\u_div/PartRem[14][2] ), .Y(\u_div/SumTmp[13][2] ) );
  MXI2X1 U159 ( .A(\u_div/SumTmp[8][2] ), .B(\u_div/PartRem[9][2] ), .S0(
        \u_div/CryTmp[8][6] ), .Y(\u_div/PartRem[8][3] ) );
  CLKINVX1 U160 ( .A(\u_div/PartRem[9][2] ), .Y(\u_div/SumTmp[8][2] ) );
  MXI2X1 U161 ( .A(\u_div/SumTmp[58][2] ), .B(\u_div/PartRem[59][2] ), .S0(
        \u_div/CryTmp[58][6] ), .Y(\u_div/PartRem[58][3] ) );
  MXI2X1 U162 ( .A(\u_div/SumTmp[57][2] ), .B(\u_div/PartRem[58][2] ), .S0(
        \u_div/CryTmp[57][6] ), .Y(\u_div/PartRem[57][3] ) );
  MXI2X1 U163 ( .A(\u_div/SumTmp[56][2] ), .B(\u_div/PartRem[57][2] ), .S0(
        \u_div/CryTmp[56][6] ), .Y(\u_div/PartRem[56][3] ) );
  MXI2X1 U164 ( .A(\u_div/SumTmp[55][2] ), .B(\u_div/PartRem[56][2] ), .S0(
        \u_div/CryTmp[55][6] ), .Y(\u_div/PartRem[55][3] ) );
  MXI2X1 U165 ( .A(\u_div/SumTmp[54][2] ), .B(\u_div/PartRem[55][2] ), .S0(
        \u_div/CryTmp[54][6] ), .Y(\u_div/PartRem[54][3] ) );
  MXI2X1 U166 ( .A(\u_div/SumTmp[52][2] ), .B(\u_div/PartRem[53][2] ), .S0(
        \u_div/CryTmp[52][6] ), .Y(\u_div/PartRem[52][3] ) );
  CLKINVX1 U167 ( .A(\u_div/PartRem[53][2] ), .Y(\u_div/SumTmp[52][2] ) );
  MXI2X1 U168 ( .A(\u_div/SumTmp[51][2] ), .B(\u_div/PartRem[52][2] ), .S0(
        \u_div/CryTmp[51][6] ), .Y(\u_div/PartRem[51][3] ) );
  CLKINVX1 U169 ( .A(\u_div/PartRem[52][2] ), .Y(\u_div/SumTmp[51][2] ) );
  MXI2X1 U170 ( .A(\u_div/SumTmp[50][2] ), .B(\u_div/PartRem[51][2] ), .S0(
        \u_div/CryTmp[50][6] ), .Y(\u_div/PartRem[50][3] ) );
  CLKINVX1 U171 ( .A(\u_div/PartRem[51][2] ), .Y(\u_div/SumTmp[50][2] ) );
  MXI2X1 U172 ( .A(\u_div/SumTmp[49][2] ), .B(\u_div/PartRem[50][2] ), .S0(
        \u_div/CryTmp[49][6] ), .Y(\u_div/PartRem[49][3] ) );
  CLKINVX1 U173 ( .A(\u_div/PartRem[50][2] ), .Y(\u_div/SumTmp[49][2] ) );
  MXI2X1 U174 ( .A(\u_div/SumTmp[47][2] ), .B(\u_div/PartRem[48][2] ), .S0(
        \u_div/CryTmp[47][6] ), .Y(\u_div/PartRem[47][3] ) );
  CLKINVX1 U175 ( .A(\u_div/PartRem[48][2] ), .Y(\u_div/SumTmp[47][2] ) );
  MXI2X1 U176 ( .A(\u_div/SumTmp[46][2] ), .B(\u_div/PartRem[47][2] ), .S0(
        \u_div/CryTmp[46][6] ), .Y(\u_div/PartRem[46][3] ) );
  CLKINVX1 U177 ( .A(\u_div/PartRem[47][2] ), .Y(\u_div/SumTmp[46][2] ) );
  MXI2X1 U178 ( .A(\u_div/SumTmp[45][2] ), .B(\u_div/PartRem[46][2] ), .S0(
        \u_div/CryTmp[45][6] ), .Y(\u_div/PartRem[45][3] ) );
  CLKINVX1 U179 ( .A(\u_div/PartRem[46][2] ), .Y(\u_div/SumTmp[45][2] ) );
  MXI2X1 U180 ( .A(\u_div/SumTmp[44][2] ), .B(\u_div/PartRem[45][2] ), .S0(
        \u_div/CryTmp[44][6] ), .Y(\u_div/PartRem[44][3] ) );
  CLKINVX1 U181 ( .A(\u_div/PartRem[45][2] ), .Y(\u_div/SumTmp[44][2] ) );
  MXI2X1 U182 ( .A(\u_div/SumTmp[42][2] ), .B(\u_div/PartRem[43][2] ), .S0(
        \u_div/CryTmp[42][6] ), .Y(\u_div/PartRem[42][3] ) );
  CLKINVX1 U183 ( .A(\u_div/PartRem[43][2] ), .Y(\u_div/SumTmp[42][2] ) );
  MXI2X1 U184 ( .A(\u_div/SumTmp[41][2] ), .B(\u_div/PartRem[42][2] ), .S0(
        \u_div/CryTmp[41][6] ), .Y(\u_div/PartRem[41][3] ) );
  CLKINVX1 U185 ( .A(\u_div/PartRem[42][2] ), .Y(\u_div/SumTmp[41][2] ) );
  MXI2X1 U186 ( .A(\u_div/SumTmp[40][2] ), .B(\u_div/PartRem[41][2] ), .S0(
        \u_div/CryTmp[40][6] ), .Y(\u_div/PartRem[40][3] ) );
  CLKINVX1 U187 ( .A(\u_div/PartRem[41][2] ), .Y(\u_div/SumTmp[40][2] ) );
  MXI2X1 U188 ( .A(\u_div/SumTmp[39][2] ), .B(\u_div/PartRem[40][2] ), .S0(
        \u_div/CryTmp[39][6] ), .Y(\u_div/PartRem[39][3] ) );
  CLKINVX1 U189 ( .A(\u_div/PartRem[40][2] ), .Y(\u_div/SumTmp[39][2] ) );
  MXI2X1 U190 ( .A(\u_div/SumTmp[37][2] ), .B(\u_div/PartRem[38][2] ), .S0(
        \u_div/CryTmp[37][6] ), .Y(\u_div/PartRem[37][3] ) );
  CLKINVX1 U191 ( .A(\u_div/PartRem[38][2] ), .Y(\u_div/SumTmp[37][2] ) );
  MXI2X1 U192 ( .A(\u_div/SumTmp[36][2] ), .B(\u_div/PartRem[37][2] ), .S0(
        \u_div/CryTmp[36][6] ), .Y(\u_div/PartRem[36][3] ) );
  CLKINVX1 U193 ( .A(\u_div/PartRem[37][2] ), .Y(\u_div/SumTmp[36][2] ) );
  MXI2X1 U194 ( .A(\u_div/SumTmp[35][2] ), .B(\u_div/PartRem[36][2] ), .S0(
        \u_div/CryTmp[35][6] ), .Y(\u_div/PartRem[35][3] ) );
  CLKINVX1 U195 ( .A(\u_div/PartRem[36][2] ), .Y(\u_div/SumTmp[35][2] ) );
  MXI2X1 U196 ( .A(\u_div/SumTmp[34][2] ), .B(\u_div/PartRem[35][2] ), .S0(
        \u_div/CryTmp[34][6] ), .Y(\u_div/PartRem[34][3] ) );
  CLKINVX1 U197 ( .A(\u_div/PartRem[35][2] ), .Y(\u_div/SumTmp[34][2] ) );
  MXI2X1 U198 ( .A(\u_div/SumTmp[32][2] ), .B(\u_div/PartRem[33][2] ), .S0(
        \u_div/CryTmp[32][6] ), .Y(\u_div/PartRem[32][3] ) );
  CLKINVX1 U199 ( .A(\u_div/PartRem[33][2] ), .Y(\u_div/SumTmp[32][2] ) );
  MXI2X1 U200 ( .A(\u_div/SumTmp[31][2] ), .B(\u_div/PartRem[32][2] ), .S0(
        \u_div/CryTmp[31][6] ), .Y(\u_div/PartRem[31][3] ) );
  CLKINVX1 U201 ( .A(\u_div/PartRem[32][2] ), .Y(\u_div/SumTmp[31][2] ) );
  MXI2X1 U202 ( .A(\u_div/SumTmp[30][2] ), .B(\u_div/PartRem[31][2] ), .S0(
        \u_div/CryTmp[30][6] ), .Y(\u_div/PartRem[30][3] ) );
  CLKINVX1 U203 ( .A(\u_div/PartRem[31][2] ), .Y(\u_div/SumTmp[30][2] ) );
  MXI2X1 U204 ( .A(\u_div/SumTmp[29][2] ), .B(\u_div/PartRem[30][2] ), .S0(
        \u_div/CryTmp[29][6] ), .Y(\u_div/PartRem[29][3] ) );
  CLKINVX1 U205 ( .A(\u_div/PartRem[30][2] ), .Y(\u_div/SumTmp[29][2] ) );
  MXI2X1 U206 ( .A(\u_div/SumTmp[27][2] ), .B(\u_div/PartRem[28][2] ), .S0(
        \u_div/CryTmp[27][6] ), .Y(\u_div/PartRem[27][3] ) );
  CLKINVX1 U207 ( .A(\u_div/PartRem[28][2] ), .Y(\u_div/SumTmp[27][2] ) );
  MXI2X1 U208 ( .A(\u_div/SumTmp[26][2] ), .B(\u_div/PartRem[27][2] ), .S0(
        \u_div/CryTmp[26][6] ), .Y(\u_div/PartRem[26][3] ) );
  CLKINVX1 U209 ( .A(\u_div/PartRem[27][2] ), .Y(\u_div/SumTmp[26][2] ) );
  MXI2X1 U210 ( .A(\u_div/SumTmp[25][2] ), .B(\u_div/PartRem[26][2] ), .S0(
        \u_div/CryTmp[25][6] ), .Y(\u_div/PartRem[25][3] ) );
  CLKINVX1 U211 ( .A(\u_div/PartRem[26][2] ), .Y(\u_div/SumTmp[25][2] ) );
  MXI2X1 U212 ( .A(\u_div/SumTmp[24][2] ), .B(\u_div/PartRem[25][2] ), .S0(
        \u_div/CryTmp[24][6] ), .Y(\u_div/PartRem[24][3] ) );
  CLKINVX1 U213 ( .A(\u_div/PartRem[25][2] ), .Y(\u_div/SumTmp[24][2] ) );
  MXI2X1 U214 ( .A(\u_div/SumTmp[22][2] ), .B(\u_div/PartRem[23][2] ), .S0(
        \u_div/CryTmp[22][6] ), .Y(\u_div/PartRem[22][3] ) );
  CLKINVX1 U215 ( .A(\u_div/PartRem[23][2] ), .Y(\u_div/SumTmp[22][2] ) );
  MXI2X1 U216 ( .A(\u_div/SumTmp[21][2] ), .B(\u_div/PartRem[22][2] ), .S0(
        \u_div/CryTmp[21][6] ), .Y(\u_div/PartRem[21][3] ) );
  CLKINVX1 U217 ( .A(\u_div/PartRem[22][2] ), .Y(\u_div/SumTmp[21][2] ) );
  MXI2X1 U218 ( .A(\u_div/SumTmp[20][2] ), .B(\u_div/PartRem[21][2] ), .S0(
        \u_div/CryTmp[20][6] ), .Y(\u_div/PartRem[20][3] ) );
  CLKINVX1 U219 ( .A(\u_div/PartRem[21][2] ), .Y(\u_div/SumTmp[20][2] ) );
  MXI2X1 U220 ( .A(\u_div/SumTmp[19][2] ), .B(\u_div/PartRem[20][2] ), .S0(
        \u_div/CryTmp[19][6] ), .Y(\u_div/PartRem[19][3] ) );
  CLKINVX1 U221 ( .A(\u_div/PartRem[20][2] ), .Y(\u_div/SumTmp[19][2] ) );
  MXI2X1 U222 ( .A(\u_div/SumTmp[17][2] ), .B(\u_div/PartRem[18][2] ), .S0(
        \u_div/CryTmp[17][6] ), .Y(\u_div/PartRem[17][3] ) );
  CLKINVX1 U223 ( .A(\u_div/PartRem[18][2] ), .Y(\u_div/SumTmp[17][2] ) );
  MXI2X1 U224 ( .A(\u_div/SumTmp[16][2] ), .B(\u_div/PartRem[17][2] ), .S0(
        \u_div/CryTmp[16][6] ), .Y(\u_div/PartRem[16][3] ) );
  CLKINVX1 U225 ( .A(\u_div/PartRem[17][2] ), .Y(\u_div/SumTmp[16][2] ) );
  MXI2X1 U226 ( .A(\u_div/SumTmp[15][2] ), .B(\u_div/PartRem[16][2] ), .S0(
        \u_div/CryTmp[15][6] ), .Y(\u_div/PartRem[15][3] ) );
  CLKINVX1 U227 ( .A(\u_div/PartRem[16][2] ), .Y(\u_div/SumTmp[15][2] ) );
  MXI2X1 U228 ( .A(\u_div/SumTmp[14][2] ), .B(\u_div/PartRem[15][2] ), .S0(
        \u_div/CryTmp[14][6] ), .Y(\u_div/PartRem[14][3] ) );
  CLKINVX1 U229 ( .A(\u_div/PartRem[15][2] ), .Y(\u_div/SumTmp[14][2] ) );
  MXI2X1 U230 ( .A(\u_div/SumTmp[12][2] ), .B(\u_div/PartRem[13][2] ), .S0(
        \u_div/CryTmp[12][6] ), .Y(\u_div/PartRem[12][3] ) );
  CLKINVX1 U231 ( .A(\u_div/PartRem[13][2] ), .Y(\u_div/SumTmp[12][2] ) );
  MXI2X1 U232 ( .A(\u_div/SumTmp[11][2] ), .B(\u_div/PartRem[12][2] ), .S0(
        \u_div/CryTmp[11][6] ), .Y(\u_div/PartRem[11][3] ) );
  CLKINVX1 U233 ( .A(\u_div/PartRem[12][2] ), .Y(\u_div/SumTmp[11][2] ) );
  MXI2X1 U234 ( .A(\u_div/SumTmp[10][2] ), .B(\u_div/PartRem[11][2] ), .S0(
        \u_div/CryTmp[10][6] ), .Y(\u_div/PartRem[10][3] ) );
  CLKINVX1 U235 ( .A(\u_div/PartRem[11][2] ), .Y(\u_div/SumTmp[10][2] ) );
  MXI2X1 U236 ( .A(\u_div/SumTmp[9][2] ), .B(\u_div/PartRem[10][2] ), .S0(
        \u_div/CryTmp[9][6] ), .Y(\u_div/PartRem[9][3] ) );
  CLKINVX1 U237 ( .A(\u_div/PartRem[10][2] ), .Y(\u_div/SumTmp[9][2] ) );
  MXI2X1 U238 ( .A(\u_div/SumTmp[7][2] ), .B(\u_div/PartRem[8][2] ), .S0(
        \u_div/CryTmp[7][6] ), .Y(\u_div/PartRem[7][3] ) );
  CLKINVX1 U239 ( .A(\u_div/PartRem[8][2] ), .Y(\u_div/SumTmp[7][2] ) );
  MXI2X1 U240 ( .A(\u_div/SumTmp[6][2] ), .B(\u_div/PartRem[7][2] ), .S0(
        \u_div/CryTmp[6][6] ), .Y(\u_div/PartRem[6][3] ) );
  CLKINVX1 U241 ( .A(\u_div/PartRem[7][2] ), .Y(\u_div/SumTmp[6][2] ) );
  MXI2X1 U242 ( .A(\u_div/SumTmp[5][2] ), .B(\u_div/PartRem[6][2] ), .S0(
        \u_div/CryTmp[5][6] ), .Y(\u_div/PartRem[5][3] ) );
  CLKINVX1 U243 ( .A(\u_div/PartRem[6][2] ), .Y(\u_div/SumTmp[5][2] ) );
  MXI2X1 U244 ( .A(\u_div/SumTmp[2][2] ), .B(\u_div/PartRem[3][2] ), .S0(
        \u_div/CryTmp[2][6] ), .Y(\u_div/PartRem[2][3] ) );
  CLKINVX1 U245 ( .A(\u_div/PartRem[3][2] ), .Y(\u_div/SumTmp[2][2] ) );
  INVX4 U246 ( .A(n2), .Y(n4) );
  INVX4 U247 ( .A(n2), .Y(n5) );
  OR2X1 U248 ( .A(\u_div/PartRem[59][5] ), .B(\u_div/u_add_PartRem_2_58/n2 ), 
        .Y(\u_div/CryTmp[58][6] ) );
  XNOR2X1 U249 ( .A(\u_div/PartRem[59][3] ), .B(\u_div/PartRem[59][2] ), .Y(
        \u_div/SumTmp[58][3] ) );
  OR2X1 U250 ( .A(\u_div/PartRem[58][5] ), .B(\u_div/u_add_PartRem_2_57/n2 ), 
        .Y(\u_div/CryTmp[57][6] ) );
  XNOR2X1 U251 ( .A(\u_div/PartRem[58][3] ), .B(\u_div/PartRem[58][2] ), .Y(
        \u_div/SumTmp[57][3] ) );
  OR2X1 U252 ( .A(\u_div/PartRem[57][5] ), .B(\u_div/u_add_PartRem_2_56/n2 ), 
        .Y(\u_div/CryTmp[56][6] ) );
  XNOR2X1 U253 ( .A(\u_div/PartRem[57][3] ), .B(\u_div/PartRem[57][2] ), .Y(
        \u_div/SumTmp[56][3] ) );
  OR2X1 U254 ( .A(\u_div/PartRem[56][5] ), .B(\u_div/u_add_PartRem_2_55/n2 ), 
        .Y(\u_div/CryTmp[55][6] ) );
  XNOR2X1 U255 ( .A(\u_div/PartRem[56][3] ), .B(\u_div/PartRem[56][2] ), .Y(
        \u_div/SumTmp[55][3] ) );
  OR2X1 U256 ( .A(\u_div/PartRem[55][5] ), .B(\u_div/u_add_PartRem_2_54/n2 ), 
        .Y(\u_div/CryTmp[54][6] ) );
  XNOR2X1 U257 ( .A(\u_div/PartRem[55][3] ), .B(\u_div/PartRem[55][2] ), .Y(
        \u_div/SumTmp[54][3] ) );
  OR2X1 U258 ( .A(\u_div/PartRem[54][5] ), .B(\u_div/u_add_PartRem_2_53/n2 ), 
        .Y(\u_div/CryTmp[53][6] ) );
  XNOR2X1 U259 ( .A(\u_div/PartRem[54][3] ), .B(\u_div/PartRem[54][2] ), .Y(
        \u_div/SumTmp[53][3] ) );
  OR2X1 U260 ( .A(\u_div/PartRem[53][5] ), .B(\u_div/u_add_PartRem_2_52/n2 ), 
        .Y(\u_div/CryTmp[52][6] ) );
  XNOR2X1 U261 ( .A(\u_div/PartRem[53][3] ), .B(\u_div/PartRem[53][2] ), .Y(
        \u_div/SumTmp[52][3] ) );
  OR2X1 U262 ( .A(\u_div/PartRem[52][5] ), .B(\u_div/u_add_PartRem_2_51/n2 ), 
        .Y(\u_div/CryTmp[51][6] ) );
  XNOR2X1 U263 ( .A(\u_div/PartRem[52][3] ), .B(\u_div/PartRem[52][2] ), .Y(
        \u_div/SumTmp[51][3] ) );
  OR2X1 U264 ( .A(\u_div/PartRem[51][5] ), .B(\u_div/u_add_PartRem_2_50/n2 ), 
        .Y(\u_div/CryTmp[50][6] ) );
  XNOR2X1 U265 ( .A(\u_div/PartRem[51][3] ), .B(\u_div/PartRem[51][2] ), .Y(
        \u_div/SumTmp[50][3] ) );
  OR2X1 U266 ( .A(\u_div/PartRem[50][5] ), .B(\u_div/u_add_PartRem_2_49/n2 ), 
        .Y(\u_div/CryTmp[49][6] ) );
  XNOR2X1 U267 ( .A(\u_div/PartRem[50][3] ), .B(\u_div/PartRem[50][2] ), .Y(
        \u_div/SumTmp[49][3] ) );
  OR2X1 U268 ( .A(\u_div/PartRem[49][5] ), .B(\u_div/u_add_PartRem_2_48/n2 ), 
        .Y(\u_div/CryTmp[48][6] ) );
  XNOR2X1 U269 ( .A(\u_div/PartRem[49][3] ), .B(\u_div/PartRem[49][2] ), .Y(
        \u_div/SumTmp[48][3] ) );
  OR2X1 U270 ( .A(\u_div/PartRem[48][5] ), .B(\u_div/u_add_PartRem_2_47/n2 ), 
        .Y(\u_div/CryTmp[47][6] ) );
  XNOR2X1 U271 ( .A(\u_div/PartRem[48][3] ), .B(\u_div/PartRem[48][2] ), .Y(
        \u_div/SumTmp[47][3] ) );
  OR2X1 U272 ( .A(\u_div/PartRem[47][5] ), .B(\u_div/u_add_PartRem_2_46/n2 ), 
        .Y(\u_div/CryTmp[46][6] ) );
  XNOR2X1 U273 ( .A(\u_div/PartRem[47][3] ), .B(\u_div/PartRem[47][2] ), .Y(
        \u_div/SumTmp[46][3] ) );
  OR2X1 U274 ( .A(\u_div/PartRem[46][5] ), .B(\u_div/u_add_PartRem_2_45/n2 ), 
        .Y(\u_div/CryTmp[45][6] ) );
  XNOR2X1 U275 ( .A(\u_div/PartRem[46][3] ), .B(\u_div/PartRem[46][2] ), .Y(
        \u_div/SumTmp[45][3] ) );
  OR2X1 U276 ( .A(\u_div/PartRem[45][5] ), .B(\u_div/u_add_PartRem_2_44/n2 ), 
        .Y(\u_div/CryTmp[44][6] ) );
  XNOR2X1 U277 ( .A(\u_div/PartRem[45][3] ), .B(\u_div/PartRem[45][2] ), .Y(
        \u_div/SumTmp[44][3] ) );
  OR2X1 U278 ( .A(\u_div/PartRem[44][5] ), .B(\u_div/u_add_PartRem_2_43/n2 ), 
        .Y(\u_div/CryTmp[43][6] ) );
  XNOR2X1 U279 ( .A(\u_div/PartRem[44][3] ), .B(\u_div/PartRem[44][2] ), .Y(
        \u_div/SumTmp[43][3] ) );
  OR2X1 U280 ( .A(\u_div/PartRem[43][5] ), .B(\u_div/u_add_PartRem_2_42/n2 ), 
        .Y(\u_div/CryTmp[42][6] ) );
  XNOR2X1 U281 ( .A(\u_div/PartRem[43][3] ), .B(\u_div/PartRem[43][2] ), .Y(
        \u_div/SumTmp[42][3] ) );
  OR2X1 U282 ( .A(\u_div/PartRem[42][5] ), .B(\u_div/u_add_PartRem_2_41/n2 ), 
        .Y(\u_div/CryTmp[41][6] ) );
  XNOR2X1 U283 ( .A(\u_div/PartRem[42][3] ), .B(\u_div/PartRem[42][2] ), .Y(
        \u_div/SumTmp[41][3] ) );
  OR2X1 U284 ( .A(\u_div/PartRem[41][5] ), .B(\u_div/u_add_PartRem_2_40/n2 ), 
        .Y(\u_div/CryTmp[40][6] ) );
  XNOR2X1 U285 ( .A(\u_div/PartRem[41][3] ), .B(\u_div/PartRem[41][2] ), .Y(
        \u_div/SumTmp[40][3] ) );
  OR2X1 U286 ( .A(\u_div/PartRem[40][5] ), .B(\u_div/u_add_PartRem_2_39/n2 ), 
        .Y(\u_div/CryTmp[39][6] ) );
  XNOR2X1 U287 ( .A(\u_div/PartRem[40][3] ), .B(\u_div/PartRem[40][2] ), .Y(
        \u_div/SumTmp[39][3] ) );
  OR2X1 U288 ( .A(\u_div/PartRem[39][5] ), .B(\u_div/u_add_PartRem_2_38/n2 ), 
        .Y(\u_div/CryTmp[38][6] ) );
  XNOR2X1 U289 ( .A(\u_div/PartRem[39][3] ), .B(\u_div/PartRem[39][2] ), .Y(
        \u_div/SumTmp[38][3] ) );
  OR2X1 U290 ( .A(\u_div/PartRem[38][5] ), .B(\u_div/u_add_PartRem_2_37/n2 ), 
        .Y(\u_div/CryTmp[37][6] ) );
  XNOR2X1 U291 ( .A(\u_div/PartRem[38][3] ), .B(\u_div/PartRem[38][2] ), .Y(
        \u_div/SumTmp[37][3] ) );
  OR2X1 U292 ( .A(\u_div/PartRem[37][5] ), .B(\u_div/u_add_PartRem_2_36/n2 ), 
        .Y(\u_div/CryTmp[36][6] ) );
  XNOR2X1 U293 ( .A(\u_div/PartRem[37][3] ), .B(\u_div/PartRem[37][2] ), .Y(
        \u_div/SumTmp[36][3] ) );
  OR2X1 U294 ( .A(\u_div/PartRem[36][5] ), .B(\u_div/u_add_PartRem_2_35/n2 ), 
        .Y(\u_div/CryTmp[35][6] ) );
  XNOR2X1 U295 ( .A(\u_div/PartRem[36][3] ), .B(\u_div/PartRem[36][2] ), .Y(
        \u_div/SumTmp[35][3] ) );
  OR2X1 U296 ( .A(\u_div/PartRem[35][5] ), .B(\u_div/u_add_PartRem_2_34/n2 ), 
        .Y(\u_div/CryTmp[34][6] ) );
  XNOR2X1 U297 ( .A(\u_div/PartRem[35][3] ), .B(\u_div/PartRem[35][2] ), .Y(
        \u_div/SumTmp[34][3] ) );
  OR2X1 U298 ( .A(\u_div/PartRem[34][5] ), .B(\u_div/u_add_PartRem_2_33/n2 ), 
        .Y(\u_div/CryTmp[33][6] ) );
  XNOR2X1 U299 ( .A(\u_div/PartRem[34][3] ), .B(\u_div/PartRem[34][2] ), .Y(
        \u_div/SumTmp[33][3] ) );
  OR2X1 U300 ( .A(\u_div/PartRem[33][5] ), .B(\u_div/u_add_PartRem_2_32/n2 ), 
        .Y(\u_div/CryTmp[32][6] ) );
  XNOR2X1 U301 ( .A(\u_div/PartRem[33][3] ), .B(\u_div/PartRem[33][2] ), .Y(
        \u_div/SumTmp[32][3] ) );
  OR2X1 U302 ( .A(\u_div/PartRem[32][5] ), .B(\u_div/u_add_PartRem_2_31/n2 ), 
        .Y(\u_div/CryTmp[31][6] ) );
  XNOR2X1 U303 ( .A(\u_div/PartRem[32][3] ), .B(\u_div/PartRem[32][2] ), .Y(
        \u_div/SumTmp[31][3] ) );
  OR2X1 U304 ( .A(\u_div/PartRem[31][5] ), .B(\u_div/u_add_PartRem_2_30/n2 ), 
        .Y(\u_div/CryTmp[30][6] ) );
  XNOR2X1 U305 ( .A(\u_div/PartRem[31][3] ), .B(\u_div/PartRem[31][2] ), .Y(
        \u_div/SumTmp[30][3] ) );
  OR2X1 U306 ( .A(\u_div/PartRem[30][5] ), .B(\u_div/u_add_PartRem_2_29/n2 ), 
        .Y(\u_div/CryTmp[29][6] ) );
  XNOR2X1 U307 ( .A(\u_div/PartRem[30][3] ), .B(\u_div/PartRem[30][2] ), .Y(
        \u_div/SumTmp[29][3] ) );
  OR2X1 U308 ( .A(\u_div/PartRem[29][5] ), .B(\u_div/u_add_PartRem_2_28/n2 ), 
        .Y(\u_div/CryTmp[28][6] ) );
  XNOR2X1 U309 ( .A(\u_div/PartRem[29][3] ), .B(\u_div/PartRem[29][2] ), .Y(
        \u_div/SumTmp[28][3] ) );
  OR2X1 U310 ( .A(\u_div/PartRem[28][5] ), .B(\u_div/u_add_PartRem_2_27/n2 ), 
        .Y(\u_div/CryTmp[27][6] ) );
  XNOR2X1 U311 ( .A(\u_div/PartRem[28][3] ), .B(\u_div/PartRem[28][2] ), .Y(
        \u_div/SumTmp[27][3] ) );
  OR2X1 U312 ( .A(\u_div/PartRem[27][5] ), .B(\u_div/u_add_PartRem_2_26/n2 ), 
        .Y(\u_div/CryTmp[26][6] ) );
  XNOR2X1 U313 ( .A(\u_div/PartRem[27][3] ), .B(\u_div/PartRem[27][2] ), .Y(
        \u_div/SumTmp[26][3] ) );
  OR2X1 U314 ( .A(\u_div/PartRem[26][5] ), .B(\u_div/u_add_PartRem_2_25/n2 ), 
        .Y(\u_div/CryTmp[25][6] ) );
  XNOR2X1 U315 ( .A(\u_div/PartRem[26][3] ), .B(\u_div/PartRem[26][2] ), .Y(
        \u_div/SumTmp[25][3] ) );
  OR2X1 U316 ( .A(\u_div/PartRem[25][5] ), .B(\u_div/u_add_PartRem_2_24/n2 ), 
        .Y(\u_div/CryTmp[24][6] ) );
  XNOR2X1 U317 ( .A(\u_div/PartRem[25][3] ), .B(\u_div/PartRem[25][2] ), .Y(
        \u_div/SumTmp[24][3] ) );
  OR2X1 U318 ( .A(\u_div/PartRem[24][5] ), .B(\u_div/u_add_PartRem_2_23/n2 ), 
        .Y(\u_div/CryTmp[23][6] ) );
  XNOR2X1 U319 ( .A(\u_div/PartRem[24][3] ), .B(\u_div/PartRem[24][2] ), .Y(
        \u_div/SumTmp[23][3] ) );
  OR2X1 U320 ( .A(\u_div/PartRem[23][5] ), .B(\u_div/u_add_PartRem_2_22/n2 ), 
        .Y(\u_div/CryTmp[22][6] ) );
  XNOR2X1 U321 ( .A(\u_div/PartRem[23][3] ), .B(\u_div/PartRem[23][2] ), .Y(
        \u_div/SumTmp[22][3] ) );
  OR2X1 U322 ( .A(\u_div/PartRem[22][5] ), .B(\u_div/u_add_PartRem_2_21/n2 ), 
        .Y(\u_div/CryTmp[21][6] ) );
  XNOR2X1 U323 ( .A(\u_div/PartRem[22][3] ), .B(\u_div/PartRem[22][2] ), .Y(
        \u_div/SumTmp[21][3] ) );
  OR2X1 U324 ( .A(\u_div/PartRem[21][5] ), .B(\u_div/u_add_PartRem_2_20/n2 ), 
        .Y(\u_div/CryTmp[20][6] ) );
  XNOR2X1 U325 ( .A(\u_div/PartRem[21][3] ), .B(\u_div/PartRem[21][2] ), .Y(
        \u_div/SumTmp[20][3] ) );
  OR2X1 U326 ( .A(\u_div/PartRem[20][5] ), .B(\u_div/u_add_PartRem_2_19/n2 ), 
        .Y(\u_div/CryTmp[19][6] ) );
  XNOR2X1 U327 ( .A(\u_div/PartRem[20][3] ), .B(\u_div/PartRem[20][2] ), .Y(
        \u_div/SumTmp[19][3] ) );
  OR2X1 U328 ( .A(\u_div/PartRem[19][5] ), .B(\u_div/u_add_PartRem_2_18/n2 ), 
        .Y(\u_div/CryTmp[18][6] ) );
  XNOR2X1 U329 ( .A(\u_div/PartRem[19][3] ), .B(\u_div/PartRem[19][2] ), .Y(
        \u_div/SumTmp[18][3] ) );
  OR2X1 U330 ( .A(\u_div/PartRem[18][5] ), .B(\u_div/u_add_PartRem_2_17/n2 ), 
        .Y(\u_div/CryTmp[17][6] ) );
  XNOR2X1 U331 ( .A(\u_div/PartRem[18][3] ), .B(\u_div/PartRem[18][2] ), .Y(
        \u_div/SumTmp[17][3] ) );
  OR2X1 U332 ( .A(\u_div/PartRem[17][5] ), .B(\u_div/u_add_PartRem_2_16/n2 ), 
        .Y(\u_div/CryTmp[16][6] ) );
  XNOR2X1 U333 ( .A(\u_div/PartRem[17][3] ), .B(\u_div/PartRem[17][2] ), .Y(
        \u_div/SumTmp[16][3] ) );
  OR2X1 U334 ( .A(\u_div/PartRem[16][5] ), .B(\u_div/u_add_PartRem_2_15/n2 ), 
        .Y(\u_div/CryTmp[15][6] ) );
  XNOR2X1 U335 ( .A(\u_div/PartRem[16][3] ), .B(\u_div/PartRem[16][2] ), .Y(
        \u_div/SumTmp[15][3] ) );
  OR2X1 U336 ( .A(\u_div/PartRem[15][5] ), .B(\u_div/u_add_PartRem_2_14/n2 ), 
        .Y(\u_div/CryTmp[14][6] ) );
  XNOR2X1 U337 ( .A(\u_div/PartRem[15][3] ), .B(\u_div/PartRem[15][2] ), .Y(
        \u_div/SumTmp[14][3] ) );
  OR2X1 U338 ( .A(\u_div/PartRem[14][5] ), .B(\u_div/u_add_PartRem_2_13/n2 ), 
        .Y(\u_div/CryTmp[13][6] ) );
  XNOR2X1 U339 ( .A(\u_div/PartRem[14][3] ), .B(\u_div/PartRem[14][2] ), .Y(
        \u_div/SumTmp[13][3] ) );
  OR2X1 U340 ( .A(\u_div/PartRem[13][5] ), .B(\u_div/u_add_PartRem_2_12/n2 ), 
        .Y(\u_div/CryTmp[12][6] ) );
  XNOR2X1 U341 ( .A(\u_div/PartRem[13][3] ), .B(\u_div/PartRem[13][2] ), .Y(
        \u_div/SumTmp[12][3] ) );
  OR2X1 U342 ( .A(\u_div/PartRem[12][5] ), .B(\u_div/u_add_PartRem_2_11/n2 ), 
        .Y(\u_div/CryTmp[11][6] ) );
  XNOR2X1 U343 ( .A(\u_div/PartRem[12][3] ), .B(\u_div/PartRem[12][2] ), .Y(
        \u_div/SumTmp[11][3] ) );
  OR2X1 U344 ( .A(\u_div/PartRem[11][5] ), .B(\u_div/u_add_PartRem_2_10/n2 ), 
        .Y(\u_div/CryTmp[10][6] ) );
  XNOR2X1 U345 ( .A(\u_div/PartRem[11][3] ), .B(\u_div/PartRem[11][2] ), .Y(
        \u_div/SumTmp[10][3] ) );
  OR2X1 U346 ( .A(\u_div/PartRem[10][5] ), .B(\u_div/u_add_PartRem_2_9/n2 ), 
        .Y(\u_div/CryTmp[9][6] ) );
  XNOR2X1 U347 ( .A(\u_div/PartRem[10][3] ), .B(\u_div/PartRem[10][2] ), .Y(
        \u_div/SumTmp[9][3] ) );
  OR2X1 U348 ( .A(\u_div/PartRem[9][5] ), .B(\u_div/u_add_PartRem_2_8/n2 ), 
        .Y(\u_div/CryTmp[8][6] ) );
  XNOR2X1 U349 ( .A(\u_div/PartRem[9][3] ), .B(\u_div/PartRem[9][2] ), .Y(
        \u_div/SumTmp[8][3] ) );
  OR2X1 U350 ( .A(\u_div/PartRem[8][5] ), .B(\u_div/u_add_PartRem_2_7/n2 ), 
        .Y(\u_div/CryTmp[7][6] ) );
  XNOR2X1 U351 ( .A(\u_div/PartRem[8][3] ), .B(\u_div/PartRem[8][2] ), .Y(
        \u_div/SumTmp[7][3] ) );
  OR2X1 U352 ( .A(\u_div/PartRem[7][5] ), .B(\u_div/u_add_PartRem_2_6/n2 ), 
        .Y(\u_div/CryTmp[6][6] ) );
  XNOR2X1 U353 ( .A(\u_div/PartRem[7][3] ), .B(\u_div/PartRem[7][2] ), .Y(
        \u_div/SumTmp[6][3] ) );
  OR2X1 U354 ( .A(\u_div/PartRem[6][5] ), .B(\u_div/u_add_PartRem_2_5/n2 ), 
        .Y(\u_div/CryTmp[5][6] ) );
  XNOR2X1 U355 ( .A(\u_div/PartRem[6][3] ), .B(\u_div/PartRem[6][2] ), .Y(
        \u_div/SumTmp[5][3] ) );
  OR2X1 U356 ( .A(\u_div/PartRem[5][5] ), .B(\u_div/u_add_PartRem_2_4/n2 ), 
        .Y(\u_div/CryTmp[4][6] ) );
  XNOR2X1 U357 ( .A(\u_div/PartRem[5][3] ), .B(\u_div/PartRem[5][2] ), .Y(
        \u_div/SumTmp[4][3] ) );
  XNOR2X1 U358 ( .A(\u_div/PartRem[4][3] ), .B(\u_div/PartRem[4][2] ), .Y(
        \u_div/SumTmp[3][3] ) );
  XNOR2X1 U359 ( .A(\u_div/PartRem[3][3] ), .B(\u_div/PartRem[3][2] ), .Y(
        \u_div/SumTmp[2][3] ) );
  XNOR2X1 U360 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/PartRem[2][2] ), .Y(
        \u_div/SumTmp[1][3] ) );
  NAND2BX1 U361 ( .AN(\u_div/PartRem[1][3] ), .B(n1), .Y(n6) );
  XNOR2X1 U362 ( .A(\u_div/PartRem[63][0] ), .B(\u_div/PartRem[62][0] ), .Y(
        \u_div/SumTmp[59][3] ) );
  XOR2X1 U363 ( .A(\u_div/CryTmp[9][6] ), .B(n3), .Y(\u_div/QInv[9] ) );
  XOR2X1 U364 ( .A(\u_div/CryTmp[8][6] ), .B(n3), .Y(\u_div/QInv[8] ) );
  XOR2X1 U365 ( .A(\u_div/CryTmp[7][6] ), .B(n4), .Y(\u_div/QInv[7] ) );
  XOR2X1 U366 ( .A(\u_div/CryTmp[6][6] ), .B(n5), .Y(\u_div/QInv[6] ) );
  XOR2X1 U367 ( .A(\u_div/CryTmp[5][6] ), .B(n4), .Y(\u_div/QInv[5] ) );
  XOR2X1 U368 ( .A(\u_div/CryTmp[59][6] ), .B(n3), .Y(\u_div/QInv[59] ) );
  XOR2X1 U369 ( .A(\u_div/CryTmp[58][6] ), .B(n5), .Y(\u_div/QInv[58] ) );
  XOR2X1 U370 ( .A(\u_div/CryTmp[57][6] ), .B(n4), .Y(\u_div/QInv[57] ) );
  XOR2X1 U371 ( .A(\u_div/CryTmp[56][6] ), .B(n3), .Y(\u_div/QInv[56] ) );
  XOR2X1 U372 ( .A(\u_div/CryTmp[55][6] ), .B(n5), .Y(\u_div/QInv[55] ) );
  XOR2X1 U373 ( .A(\u_div/CryTmp[54][6] ), .B(n4), .Y(\u_div/QInv[54] ) );
  XOR2X1 U374 ( .A(\u_div/CryTmp[53][6] ), .B(n3), .Y(\u_div/QInv[53] ) );
  XOR2X1 U375 ( .A(\u_div/CryTmp[50][6] ), .B(n3), .Y(\u_div/QInv[50] ) );
  XOR2X1 U376 ( .A(\u_div/CryTmp[4][6] ), .B(n5), .Y(\u_div/QInv[4] ) );
  XOR2X1 U377 ( .A(\u_div/CryTmp[49][6] ), .B(n4), .Y(\u_div/QInv[49] ) );
  XOR2X1 U378 ( .A(\u_div/CryTmp[48][6] ), .B(n3), .Y(\u_div/QInv[48] ) );
  XOR2X1 U379 ( .A(\u_div/CryTmp[47][6] ), .B(n5), .Y(\u_div/QInv[47] ) );
  XOR2X1 U380 ( .A(\u_div/CryTmp[46][6] ), .B(n4), .Y(\u_div/QInv[46] ) );
  XOR2X1 U381 ( .A(\u_div/CryTmp[45][6] ), .B(n3), .Y(\u_div/QInv[45] ) );
  XOR2X1 U382 ( .A(\u_div/CryTmp[44][6] ), .B(n5), .Y(\u_div/QInv[44] ) );
  XOR2X1 U383 ( .A(\u_div/CryTmp[43][6] ), .B(n4), .Y(\u_div/QInv[43] ) );
  XOR2X1 U384 ( .A(\u_div/CryTmp[42][6] ), .B(n3), .Y(\u_div/QInv[42] ) );
  XOR2X1 U385 ( .A(\u_div/CryTmp[40][6] ), .B(n4), .Y(\u_div/QInv[40] ) );
  XOR2X1 U386 ( .A(\u_div/CryTmp[39][6] ), .B(n5), .Y(\u_div/QInv[39] ) );
  XOR2X1 U387 ( .A(\u_div/CryTmp[38][6] ), .B(n4), .Y(\u_div/QInv[38] ) );
  XOR2X1 U388 ( .A(\u_div/CryTmp[37][6] ), .B(n3), .Y(\u_div/QInv[37] ) );
  XOR2X1 U389 ( .A(\u_div/CryTmp[36][6] ), .B(n5), .Y(\u_div/QInv[36] ) );
  XOR2X1 U390 ( .A(\u_div/CryTmp[35][6] ), .B(n4), .Y(\u_div/QInv[35] ) );
  XOR2X1 U391 ( .A(\u_div/CryTmp[34][6] ), .B(n5), .Y(\u_div/QInv[34] ) );
  XOR2X1 U392 ( .A(\u_div/CryTmp[33][6] ), .B(n4), .Y(\u_div/QInv[33] ) );
  XOR2X1 U393 ( .A(\u_div/CryTmp[30][6] ), .B(n4), .Y(\u_div/QInv[30] ) );
  XOR2X1 U394 ( .A(\u_div/CryTmp[2][6] ), .B(n3), .Y(\u_div/QInv[2] ) );
  XOR2X1 U395 ( .A(\u_div/CryTmp[29][6] ), .B(n5), .Y(\u_div/QInv[29] ) );
  XOR2X1 U396 ( .A(\u_div/CryTmp[28][6] ), .B(n4), .Y(\u_div/QInv[28] ) );
  XOR2X1 U397 ( .A(\u_div/CryTmp[27][6] ), .B(n3), .Y(\u_div/QInv[27] ) );
  XOR2X1 U398 ( .A(\u_div/CryTmp[26][6] ), .B(n5), .Y(\u_div/QInv[26] ) );
  XOR2X1 U399 ( .A(\u_div/CryTmp[25][6] ), .B(n4), .Y(\u_div/QInv[25] ) );
  XOR2X1 U400 ( .A(\u_div/CryTmp[24][6] ), .B(n3), .Y(\u_div/QInv[24] ) );
  XOR2X1 U401 ( .A(\u_div/CryTmp[23][6] ), .B(n5), .Y(\u_div/QInv[23] ) );
  XOR2X1 U402 ( .A(\u_div/CryTmp[20][6] ), .B(n5), .Y(\u_div/QInv[20] ) );
  XOR2X1 U403 ( .A(\u_div/CryTmp[19][6] ), .B(n3), .Y(\u_div/QInv[19] ) );
  XOR2X1 U404 ( .A(\u_div/CryTmp[18][6] ), .B(n5), .Y(\u_div/QInv[18] ) );
  XOR2X1 U405 ( .A(\u_div/CryTmp[17][6] ), .B(n4), .Y(\u_div/QInv[17] ) );
  XOR2X1 U406 ( .A(\u_div/CryTmp[16][6] ), .B(n5), .Y(\u_div/QInv[16] ) );
  XOR2X1 U407 ( .A(\u_div/CryTmp[15][6] ), .B(n4), .Y(\u_div/QInv[15] ) );
  XOR2X1 U408 ( .A(\u_div/CryTmp[14][6] ), .B(n5), .Y(\u_div/QInv[14] ) );
  XOR2X1 U409 ( .A(\u_div/CryTmp[13][6] ), .B(n4), .Y(\u_div/QInv[13] ) );
  XOR2X1 U410 ( .A(\u_div/CryTmp[10][6] ), .B(n5), .Y(\u_div/QInv[10] ) );
endmodule


module GSIM_DW01_inc_4 ( A, SUM );
  input [63:0] A;
  output [63:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;

  NOR3BX1 U2 ( .AN(A[59]), .B(n1), .C(n24), .Y(n22) );
  NOR3BX1 U3 ( .AN(A[55]), .B(n2), .C(n30), .Y(n28) );
  NOR3BX1 U4 ( .AN(A[51]), .B(n3), .C(n34), .Y(n32) );
  NOR3BX1 U5 ( .AN(A[47]), .B(n4), .C(n38), .Y(n36) );
  NOR3BX1 U6 ( .AN(A[43]), .B(n5), .C(n42), .Y(n40) );
  NOR3BX1 U7 ( .AN(A[39]), .B(n6), .C(n46), .Y(n44) );
  NOR3BX1 U8 ( .AN(A[35]), .B(n7), .C(n52), .Y(n50) );
  NOR3BX1 U9 ( .AN(A[31]), .B(n8), .C(n56), .Y(n54) );
  NOR3BX1 U10 ( .AN(A[27]), .B(n9), .C(n60), .Y(n58) );
  NOR3BX1 U11 ( .AN(A[23]), .B(n10), .C(n64), .Y(n62) );
  NOR3BX1 U12 ( .AN(A[19]), .B(n11), .C(n68), .Y(n66) );
  NOR3BX1 U13 ( .AN(A[15]), .B(n12), .C(n72), .Y(n70) );
  NOR3BX1 U14 ( .AN(A[11]), .B(n13), .C(n76), .Y(n74) );
  NOR3BX1 U15 ( .AN(A[7]), .B(n14), .C(n19), .Y(n17) );
  NAND3X1 U16 ( .A(A[4]), .B(n26), .C(A[5]), .Y(n19) );
  NAND2X1 U17 ( .A(A[60]), .B(n22), .Y(n23) );
  NOR3BX1 U18 ( .AN(A[3]), .B(n15), .C(n48), .Y(n26) );
  NOR2XL U19 ( .A(n24), .B(n1), .Y(n27) );
  NAND2XL U20 ( .A(A[56]), .B(n28), .Y(n29) );
  NOR2XL U21 ( .A(n30), .B(n2), .Y(n31) );
  NAND2XL U22 ( .A(A[52]), .B(n32), .Y(n33) );
  NOR2XL U23 ( .A(n34), .B(n3), .Y(n35) );
  NAND2XL U24 ( .A(A[48]), .B(n36), .Y(n37) );
  NOR2XL U25 ( .A(n38), .B(n4), .Y(n39) );
  NAND2XL U26 ( .A(A[44]), .B(n40), .Y(n41) );
  NOR2XL U27 ( .A(n42), .B(n5), .Y(n43) );
  NAND2XL U28 ( .A(A[40]), .B(n44), .Y(n45) );
  NOR2XL U29 ( .A(n46), .B(n6), .Y(n49) );
  NAND2XL U30 ( .A(A[36]), .B(n50), .Y(n51) );
  NOR2XL U31 ( .A(n52), .B(n7), .Y(n53) );
  NAND2XL U32 ( .A(A[32]), .B(n54), .Y(n55) );
  NOR2XL U33 ( .A(n56), .B(n8), .Y(n57) );
  NAND2XL U34 ( .A(A[28]), .B(n58), .Y(n59) );
  NOR2XL U35 ( .A(n60), .B(n9), .Y(n61) );
  NAND2XL U36 ( .A(A[24]), .B(n62), .Y(n63) );
  NOR2XL U37 ( .A(n64), .B(n10), .Y(n65) );
  NAND2XL U38 ( .A(A[20]), .B(n66), .Y(n67) );
  NOR2XL U39 ( .A(n68), .B(n11), .Y(n69) );
  NAND2XL U40 ( .A(A[16]), .B(n70), .Y(n71) );
  NOR2XL U41 ( .A(n72), .B(n12), .Y(n73) );
  NAND2XL U42 ( .A(A[12]), .B(n74), .Y(n75) );
  NOR2XL U43 ( .A(n76), .B(n13), .Y(n77) );
  NAND2XL U44 ( .A(A[8]), .B(n17), .Y(n16) );
  NOR2XL U45 ( .A(n19), .B(n14), .Y(n18) );
  NAND2XL U46 ( .A(A[4]), .B(n26), .Y(n25) );
  XNOR2XL U47 ( .A(A[61]), .B(n23), .Y(SUM[61]) );
  XOR2XL U48 ( .A(A[60]), .B(n22), .Y(SUM[60]) );
  XNOR2XL U49 ( .A(A[62]), .B(n21), .Y(SUM[62]) );
  NOR2XL U50 ( .A(n48), .B(n15), .Y(n47) );
  CLKINVX1 U51 ( .A(A[58]), .Y(n1) );
  CLKINVX1 U52 ( .A(A[54]), .Y(n2) );
  CLKINVX1 U53 ( .A(A[50]), .Y(n3) );
  CLKINVX1 U54 ( .A(A[46]), .Y(n4) );
  CLKINVX1 U55 ( .A(A[42]), .Y(n5) );
  CLKINVX1 U56 ( .A(A[38]), .Y(n6) );
  CLKINVX1 U57 ( .A(A[34]), .Y(n7) );
  CLKINVX1 U58 ( .A(A[30]), .Y(n8) );
  CLKINVX1 U59 ( .A(A[26]), .Y(n9) );
  CLKINVX1 U60 ( .A(A[22]), .Y(n10) );
  CLKINVX1 U61 ( .A(A[2]), .Y(n15) );
  CLKINVX1 U62 ( .A(A[18]), .Y(n11) );
  CLKINVX1 U63 ( .A(A[6]), .Y(n14) );
  CLKINVX1 U64 ( .A(A[14]), .Y(n12) );
  CLKINVX1 U65 ( .A(A[10]), .Y(n13) );
  XNOR2X1 U66 ( .A(A[9]), .B(n16), .Y(SUM[9]) );
  XOR2X1 U67 ( .A(A[8]), .B(n17), .Y(SUM[8]) );
  XOR2X1 U68 ( .A(A[7]), .B(n18), .Y(SUM[7]) );
  XOR2X1 U69 ( .A(n14), .B(n19), .Y(SUM[6]) );
  XOR2X1 U70 ( .A(A[63]), .B(n20), .Y(SUM[63]) );
  NOR2BX1 U71 ( .AN(A[62]), .B(n21), .Y(n20) );
  NAND3X1 U72 ( .A(A[60]), .B(n22), .C(A[61]), .Y(n21) );
  XNOR2X1 U73 ( .A(A[5]), .B(n25), .Y(SUM[5]) );
  XOR2X1 U74 ( .A(A[59]), .B(n27), .Y(SUM[59]) );
  XOR2X1 U75 ( .A(n1), .B(n24), .Y(SUM[58]) );
  NAND3X1 U76 ( .A(A[56]), .B(n28), .C(A[57]), .Y(n24) );
  XNOR2X1 U77 ( .A(A[57]), .B(n29), .Y(SUM[57]) );
  XOR2X1 U78 ( .A(A[56]), .B(n28), .Y(SUM[56]) );
  XOR2X1 U79 ( .A(A[55]), .B(n31), .Y(SUM[55]) );
  XOR2X1 U80 ( .A(n2), .B(n30), .Y(SUM[54]) );
  NAND3X1 U81 ( .A(A[52]), .B(n32), .C(A[53]), .Y(n30) );
  XNOR2X1 U82 ( .A(A[53]), .B(n33), .Y(SUM[53]) );
  XOR2X1 U83 ( .A(A[52]), .B(n32), .Y(SUM[52]) );
  XOR2X1 U84 ( .A(A[51]), .B(n35), .Y(SUM[51]) );
  XOR2X1 U85 ( .A(n3), .B(n34), .Y(SUM[50]) );
  NAND3X1 U86 ( .A(A[48]), .B(n36), .C(A[49]), .Y(n34) );
  XOR2X1 U87 ( .A(A[4]), .B(n26), .Y(SUM[4]) );
  XNOR2X1 U88 ( .A(A[49]), .B(n37), .Y(SUM[49]) );
  XOR2X1 U89 ( .A(A[48]), .B(n36), .Y(SUM[48]) );
  XOR2X1 U90 ( .A(A[47]), .B(n39), .Y(SUM[47]) );
  XOR2X1 U91 ( .A(n4), .B(n38), .Y(SUM[46]) );
  NAND3X1 U92 ( .A(A[44]), .B(n40), .C(A[45]), .Y(n38) );
  XNOR2X1 U93 ( .A(A[45]), .B(n41), .Y(SUM[45]) );
  XOR2X1 U94 ( .A(A[44]), .B(n40), .Y(SUM[44]) );
  XOR2X1 U95 ( .A(A[43]), .B(n43), .Y(SUM[43]) );
  XOR2X1 U96 ( .A(n5), .B(n42), .Y(SUM[42]) );
  NAND3X1 U97 ( .A(A[40]), .B(n44), .C(A[41]), .Y(n42) );
  XNOR2X1 U98 ( .A(A[41]), .B(n45), .Y(SUM[41]) );
  XOR2X1 U99 ( .A(A[40]), .B(n44), .Y(SUM[40]) );
  XOR2X1 U100 ( .A(A[3]), .B(n47), .Y(SUM[3]) );
  XOR2X1 U101 ( .A(A[39]), .B(n49), .Y(SUM[39]) );
  XOR2X1 U102 ( .A(n6), .B(n46), .Y(SUM[38]) );
  NAND3X1 U103 ( .A(A[36]), .B(n50), .C(A[37]), .Y(n46) );
  XNOR2X1 U104 ( .A(A[37]), .B(n51), .Y(SUM[37]) );
  XOR2X1 U105 ( .A(A[36]), .B(n50), .Y(SUM[36]) );
  XOR2X1 U106 ( .A(A[35]), .B(n53), .Y(SUM[35]) );
  XOR2X1 U107 ( .A(n7), .B(n52), .Y(SUM[34]) );
  NAND3X1 U108 ( .A(A[32]), .B(n54), .C(A[33]), .Y(n52) );
  XNOR2X1 U109 ( .A(A[33]), .B(n55), .Y(SUM[33]) );
  XOR2X1 U110 ( .A(A[32]), .B(n54), .Y(SUM[32]) );
  XOR2X1 U111 ( .A(A[31]), .B(n57), .Y(SUM[31]) );
  XOR2X1 U112 ( .A(n8), .B(n56), .Y(SUM[30]) );
  NAND3X1 U113 ( .A(A[28]), .B(n58), .C(A[29]), .Y(n56) );
  XOR2X1 U114 ( .A(n15), .B(n48), .Y(SUM[2]) );
  XNOR2X1 U115 ( .A(A[29]), .B(n59), .Y(SUM[29]) );
  XOR2X1 U116 ( .A(A[28]), .B(n58), .Y(SUM[28]) );
  XOR2X1 U117 ( .A(A[27]), .B(n61), .Y(SUM[27]) );
  XOR2X1 U118 ( .A(n9), .B(n60), .Y(SUM[26]) );
  NAND3X1 U119 ( .A(A[24]), .B(n62), .C(A[25]), .Y(n60) );
  XNOR2X1 U120 ( .A(A[25]), .B(n63), .Y(SUM[25]) );
  XOR2X1 U121 ( .A(A[24]), .B(n62), .Y(SUM[24]) );
  XOR2X1 U122 ( .A(A[23]), .B(n65), .Y(SUM[23]) );
  XOR2X1 U123 ( .A(n10), .B(n64), .Y(SUM[22]) );
  NAND3X1 U124 ( .A(A[20]), .B(n66), .C(A[21]), .Y(n64) );
  XNOR2X1 U125 ( .A(A[21]), .B(n67), .Y(SUM[21]) );
  XOR2X1 U126 ( .A(A[20]), .B(n66), .Y(SUM[20]) );
  XOR2X1 U127 ( .A(A[19]), .B(n69), .Y(SUM[19]) );
  XOR2X1 U128 ( .A(n11), .B(n68), .Y(SUM[18]) );
  NAND3X1 U129 ( .A(A[16]), .B(n70), .C(A[17]), .Y(n68) );
  XNOR2X1 U130 ( .A(A[17]), .B(n71), .Y(SUM[17]) );
  XOR2X1 U131 ( .A(A[16]), .B(n70), .Y(SUM[16]) );
  XOR2X1 U132 ( .A(A[15]), .B(n73), .Y(SUM[15]) );
  XOR2X1 U133 ( .A(n12), .B(n72), .Y(SUM[14]) );
  NAND3X1 U134 ( .A(A[12]), .B(n74), .C(A[13]), .Y(n72) );
  XNOR2X1 U135 ( .A(A[13]), .B(n75), .Y(SUM[13]) );
  XOR2X1 U136 ( .A(A[12]), .B(n74), .Y(SUM[12]) );
  XOR2X1 U137 ( .A(A[11]), .B(n77), .Y(SUM[11]) );
  XOR2X1 U138 ( .A(n13), .B(n76), .Y(SUM[10]) );
  NAND3X1 U139 ( .A(A[8]), .B(n17), .C(A[9]), .Y(n76) );
  NAND2X1 U140 ( .A(A[1]), .B(A[0]), .Y(n48) );
endmodule


module GSIM_DW01_absval_2 ( A, ABSVAL );
  input [63:0] A;
  output [63:0] ABSVAL;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68;
  wire   [63:0] AMUX1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  GSIM_DW01_inc_4 NEG ( .A({n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
        n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
        n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
        n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
        n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68}), .SUM({
        AMUX1[63:2], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1}) );
  INVX1 U1 ( .A(A[63]), .Y(n5) );
  CLKMX2X2 U2 ( .A(A[61]), .B(AMUX1[61]), .S0(n4), .Y(ABSVAL[61]) );
  CLKINVX1 U3 ( .A(A[61]), .Y(n7) );
  INVX3 U4 ( .A(n5), .Y(n4) );
  INVX3 U5 ( .A(n5), .Y(n3) );
  INVX3 U6 ( .A(n5), .Y(n2) );
  INVX3 U7 ( .A(n5), .Y(n1) );
  CLKINVX1 U8 ( .A(A[59]), .Y(n9) );
  CLKINVX1 U9 ( .A(A[60]), .Y(n8) );
  CLKINVX1 U10 ( .A(A[58]), .Y(n10) );
  CLKINVX1 U11 ( .A(A[54]), .Y(n14) );
  CLKINVX1 U12 ( .A(A[50]), .Y(n18) );
  CLKINVX1 U13 ( .A(A[46]), .Y(n22) );
  CLKINVX1 U14 ( .A(A[42]), .Y(n26) );
  CLKINVX1 U15 ( .A(A[57]), .Y(n11) );
  CLKINVX1 U16 ( .A(A[53]), .Y(n15) );
  CLKINVX1 U17 ( .A(A[49]), .Y(n19) );
  CLKINVX1 U18 ( .A(A[62]), .Y(n6) );
  CLKINVX1 U19 ( .A(A[55]), .Y(n13) );
  CLKINVX1 U20 ( .A(A[51]), .Y(n17) );
  CLKINVX1 U21 ( .A(A[47]), .Y(n21) );
  CLKINVX1 U22 ( .A(A[43]), .Y(n25) );
  CLKINVX1 U23 ( .A(A[39]), .Y(n29) );
  CLKINVX1 U24 ( .A(A[35]), .Y(n33) );
  CLKINVX1 U25 ( .A(A[31]), .Y(n37) );
  CLKINVX1 U26 ( .A(A[56]), .Y(n12) );
  CLKINVX1 U27 ( .A(A[52]), .Y(n16) );
  CLKINVX1 U28 ( .A(A[48]), .Y(n20) );
  CLKINVX1 U29 ( .A(A[44]), .Y(n24) );
  CLKINVX1 U30 ( .A(A[40]), .Y(n28) );
  CLKINVX1 U31 ( .A(A[36]), .Y(n32) );
  CLKINVX1 U32 ( .A(A[32]), .Y(n36) );
  CLKINVX1 U33 ( .A(A[38]), .Y(n30) );
  CLKINVX1 U34 ( .A(A[34]), .Y(n34) );
  CLKINVX1 U35 ( .A(A[30]), .Y(n38) );
  CLKINVX1 U36 ( .A(A[26]), .Y(n42) );
  CLKINVX1 U37 ( .A(A[22]), .Y(n46) );
  CLKINVX1 U38 ( .A(A[2]), .Y(n66) );
  CLKINVX1 U39 ( .A(A[45]), .Y(n23) );
  CLKINVX1 U40 ( .A(A[41]), .Y(n27) );
  CLKINVX1 U41 ( .A(A[37]), .Y(n31) );
  CLKINVX1 U42 ( .A(A[33]), .Y(n35) );
  CLKINVX1 U43 ( .A(A[29]), .Y(n39) );
  CLKINVX1 U44 ( .A(A[25]), .Y(n43) );
  CLKINVX1 U45 ( .A(A[21]), .Y(n47) );
  CLKINVX1 U46 ( .A(A[27]), .Y(n41) );
  CLKINVX1 U47 ( .A(A[23]), .Y(n45) );
  CLKINVX1 U48 ( .A(A[19]), .Y(n49) );
  CLKINVX1 U49 ( .A(A[15]), .Y(n53) );
  CLKINVX1 U50 ( .A(A[11]), .Y(n57) );
  CLKINVX1 U51 ( .A(A[7]), .Y(n61) );
  CLKINVX1 U52 ( .A(A[3]), .Y(n65) );
  CLKINVX1 U53 ( .A(A[18]), .Y(n50) );
  CLKINVX1 U54 ( .A(A[28]), .Y(n40) );
  CLKINVX1 U55 ( .A(A[24]), .Y(n44) );
  CLKINVX1 U56 ( .A(A[20]), .Y(n48) );
  CLKINVX1 U57 ( .A(A[16]), .Y(n52) );
  CLKINVX1 U58 ( .A(A[12]), .Y(n56) );
  CLKINVX1 U59 ( .A(A[8]), .Y(n60) );
  CLKINVX1 U60 ( .A(A[4]), .Y(n64) );
  CLKINVX1 U61 ( .A(A[6]), .Y(n62) );
  CLKINVX1 U62 ( .A(A[17]), .Y(n51) );
  CLKINVX1 U63 ( .A(A[13]), .Y(n55) );
  CLKINVX1 U64 ( .A(A[9]), .Y(n59) );
  CLKINVX1 U65 ( .A(A[5]), .Y(n63) );
  CLKINVX1 U66 ( .A(A[14]), .Y(n54) );
  CLKINVX1 U67 ( .A(A[10]), .Y(n58) );
  CLKINVX1 U68 ( .A(A[0]), .Y(n68) );
  CLKINVX1 U69 ( .A(A[1]), .Y(n67) );
  CLKMX2X2 U70 ( .A(A[9]), .B(AMUX1[9]), .S0(n3), .Y(ABSVAL[9]) );
  CLKMX2X2 U71 ( .A(A[8]), .B(AMUX1[8]), .S0(n4), .Y(ABSVAL[8]) );
  CLKMX2X2 U72 ( .A(A[7]), .B(AMUX1[7]), .S0(n4), .Y(ABSVAL[7]) );
  CLKMX2X2 U73 ( .A(A[6]), .B(AMUX1[6]), .S0(n4), .Y(ABSVAL[6]) );
  AND2X1 U74 ( .A(AMUX1[63]), .B(n4), .Y(ABSVAL[63]) );
  CLKMX2X2 U75 ( .A(A[62]), .B(AMUX1[62]), .S0(n4), .Y(ABSVAL[62]) );
  CLKMX2X2 U76 ( .A(A[60]), .B(AMUX1[60]), .S0(n4), .Y(ABSVAL[60]) );
  CLKMX2X2 U77 ( .A(A[5]), .B(AMUX1[5]), .S0(n4), .Y(ABSVAL[5]) );
  CLKMX2X2 U78 ( .A(A[59]), .B(AMUX1[59]), .S0(n4), .Y(ABSVAL[59]) );
  CLKMX2X2 U79 ( .A(A[58]), .B(AMUX1[58]), .S0(n4), .Y(ABSVAL[58]) );
  CLKMX2X2 U80 ( .A(A[57]), .B(AMUX1[57]), .S0(n4), .Y(ABSVAL[57]) );
  CLKMX2X2 U81 ( .A(A[56]), .B(AMUX1[56]), .S0(n3), .Y(ABSVAL[56]) );
  CLKMX2X2 U82 ( .A(A[55]), .B(AMUX1[55]), .S0(n3), .Y(ABSVAL[55]) );
  CLKMX2X2 U83 ( .A(A[54]), .B(AMUX1[54]), .S0(n3), .Y(ABSVAL[54]) );
  CLKMX2X2 U84 ( .A(A[53]), .B(AMUX1[53]), .S0(n3), .Y(ABSVAL[53]) );
  CLKMX2X2 U85 ( .A(A[52]), .B(AMUX1[52]), .S0(n3), .Y(ABSVAL[52]) );
  CLKMX2X2 U86 ( .A(A[51]), .B(AMUX1[51]), .S0(n3), .Y(ABSVAL[51]) );
  CLKMX2X2 U87 ( .A(A[50]), .B(AMUX1[50]), .S0(n3), .Y(ABSVAL[50]) );
  CLKMX2X2 U88 ( .A(A[4]), .B(AMUX1[4]), .S0(n3), .Y(ABSVAL[4]) );
  CLKMX2X2 U89 ( .A(A[49]), .B(AMUX1[49]), .S0(n3), .Y(ABSVAL[49]) );
  CLKMX2X2 U90 ( .A(A[48]), .B(AMUX1[48]), .S0(n3), .Y(ABSVAL[48]) );
  CLKMX2X2 U91 ( .A(A[47]), .B(AMUX1[47]), .S0(n3), .Y(ABSVAL[47]) );
  CLKMX2X2 U92 ( .A(A[46]), .B(AMUX1[46]), .S0(n3), .Y(ABSVAL[46]) );
  CLKMX2X2 U93 ( .A(A[45]), .B(AMUX1[45]), .S0(n3), .Y(ABSVAL[45]) );
  CLKMX2X2 U94 ( .A(A[44]), .B(AMUX1[44]), .S0(n2), .Y(ABSVAL[44]) );
  CLKMX2X2 U95 ( .A(A[43]), .B(AMUX1[43]), .S0(n2), .Y(ABSVAL[43]) );
  CLKMX2X2 U96 ( .A(A[42]), .B(AMUX1[42]), .S0(n2), .Y(ABSVAL[42]) );
  CLKMX2X2 U97 ( .A(A[41]), .B(AMUX1[41]), .S0(n2), .Y(ABSVAL[41]) );
  CLKMX2X2 U98 ( .A(A[40]), .B(AMUX1[40]), .S0(n2), .Y(ABSVAL[40]) );
  CLKMX2X2 U99 ( .A(A[3]), .B(AMUX1[3]), .S0(n2), .Y(ABSVAL[3]) );
  CLKMX2X2 U100 ( .A(A[39]), .B(AMUX1[39]), .S0(n2), .Y(ABSVAL[39]) );
  CLKMX2X2 U101 ( .A(A[38]), .B(AMUX1[38]), .S0(n2), .Y(ABSVAL[38]) );
  CLKMX2X2 U102 ( .A(A[37]), .B(AMUX1[37]), .S0(n2), .Y(ABSVAL[37]) );
  CLKMX2X2 U103 ( .A(A[36]), .B(AMUX1[36]), .S0(n2), .Y(ABSVAL[36]) );
  CLKMX2X2 U104 ( .A(A[35]), .B(AMUX1[35]), .S0(n2), .Y(ABSVAL[35]) );
  CLKMX2X2 U105 ( .A(A[34]), .B(AMUX1[34]), .S0(n2), .Y(ABSVAL[34]) );
  CLKMX2X2 U106 ( .A(A[33]), .B(AMUX1[33]), .S0(n1), .Y(ABSVAL[33]) );
  CLKMX2X2 U107 ( .A(A[32]), .B(AMUX1[32]), .S0(n1), .Y(ABSVAL[32]) );
  CLKMX2X2 U108 ( .A(A[31]), .B(AMUX1[31]), .S0(n1), .Y(ABSVAL[31]) );
  CLKMX2X2 U109 ( .A(A[30]), .B(AMUX1[30]), .S0(n1), .Y(ABSVAL[30]) );
  CLKMX2X2 U110 ( .A(A[2]), .B(AMUX1[2]), .S0(n1), .Y(ABSVAL[2]) );
  CLKMX2X2 U111 ( .A(A[29]), .B(AMUX1[29]), .S0(n1), .Y(ABSVAL[29]) );
  CLKMX2X2 U112 ( .A(A[28]), .B(AMUX1[28]), .S0(n1), .Y(ABSVAL[28]) );
  CLKMX2X2 U113 ( .A(A[27]), .B(AMUX1[27]), .S0(n1), .Y(ABSVAL[27]) );
  CLKMX2X2 U114 ( .A(A[26]), .B(AMUX1[26]), .S0(n1), .Y(ABSVAL[26]) );
  CLKMX2X2 U115 ( .A(A[25]), .B(AMUX1[25]), .S0(n1), .Y(ABSVAL[25]) );
  CLKMX2X2 U116 ( .A(A[24]), .B(AMUX1[24]), .S0(n1), .Y(ABSVAL[24]) );
  CLKMX2X2 U117 ( .A(A[23]), .B(AMUX1[23]), .S0(n1), .Y(ABSVAL[23]) );
  CLKMX2X2 U118 ( .A(A[22]), .B(AMUX1[22]), .S0(n1), .Y(ABSVAL[22]) );
  CLKMX2X2 U119 ( .A(A[21]), .B(AMUX1[21]), .S0(n1), .Y(ABSVAL[21]) );
  CLKMX2X2 U120 ( .A(A[20]), .B(AMUX1[20]), .S0(n1), .Y(ABSVAL[20]) );
  CLKMX2X2 U121 ( .A(A[19]), .B(AMUX1[19]), .S0(n1), .Y(ABSVAL[19]) );
  CLKMX2X2 U122 ( .A(A[18]), .B(AMUX1[18]), .S0(n1), .Y(ABSVAL[18]) );
  CLKMX2X2 U123 ( .A(A[17]), .B(AMUX1[17]), .S0(n2), .Y(ABSVAL[17]) );
  CLKMX2X2 U124 ( .A(A[16]), .B(AMUX1[16]), .S0(n2), .Y(ABSVAL[16]) );
  CLKMX2X2 U125 ( .A(A[15]), .B(AMUX1[15]), .S0(n2), .Y(ABSVAL[15]) );
  CLKMX2X2 U126 ( .A(A[14]), .B(AMUX1[14]), .S0(n2), .Y(ABSVAL[14]) );
  CLKMX2X2 U127 ( .A(A[13]), .B(AMUX1[13]), .S0(n3), .Y(ABSVAL[13]) );
  CLKMX2X2 U128 ( .A(A[12]), .B(AMUX1[12]), .S0(n3), .Y(ABSVAL[12]) );
  CLKMX2X2 U129 ( .A(A[11]), .B(AMUX1[11]), .S0(n3), .Y(ABSVAL[11]) );
  CLKMX2X2 U130 ( .A(A[10]), .B(AMUX1[10]), .S0(n2), .Y(ABSVAL[10]) );
endmodule


module GSIM_DW_inc_2 ( carry_in, a, carry_out, sum );
  input [63:0] a;
  output [63:0] sum;
  input carry_in;
  output carry_out;
  wire   \sum[63] , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63;
  assign sum[62] = \sum[63] ;
  assign sum[61] = \sum[63] ;
  assign sum[63] = \sum[63] ;

  ADDHXL U8 ( .A(a[58]), .B(n6), .CO(n5), .S(sum[58]) );
  ADDHXL U10 ( .A(a[56]), .B(n8), .CO(n7), .S(sum[56]) );
  ADDHXL U13 ( .A(a[53]), .B(n11), .CO(n10), .S(sum[53]) );
  ADDHXL U16 ( .A(a[50]), .B(n14), .CO(n13), .S(sum[50]) );
  ADDHXL U18 ( .A(a[48]), .B(n16), .CO(n15), .S(sum[48]) );
  ADDHXL U21 ( .A(a[45]), .B(n19), .CO(n18), .S(sum[45]) );
  ADDHXL U24 ( .A(a[42]), .B(n22), .CO(n21), .S(sum[42]) );
  ADDHXL U27 ( .A(a[39]), .B(n25), .CO(n24), .S(sum[39]) );
  ADDHXL U29 ( .A(a[37]), .B(n27), .CO(n26), .S(sum[37]) );
  ADDHXL U32 ( .A(a[34]), .B(n30), .CO(n29), .S(sum[34]) );
  ADDHXL U36 ( .A(a[30]), .B(n34), .CO(n33), .S(sum[30]) );
  ADDHXL U39 ( .A(a[27]), .B(n37), .CO(n36), .S(sum[27]) );
  ADDHXL U42 ( .A(a[24]), .B(n40), .CO(n39), .S(sum[24]) );
  ADDHXL U45 ( .A(a[21]), .B(n43), .CO(n42), .S(sum[21]) );
  ADDHXL U47 ( .A(a[19]), .B(n45), .CO(n44), .S(sum[19]) );
  ADDHXL U54 ( .A(a[12]), .B(n52), .CO(n51), .S(sum[12]) );
  ADDHXL U55 ( .A(a[11]), .B(n53), .CO(n52), .S(sum[11]) );
  ADDHXL U57 ( .A(a[9]), .B(n55), .CO(n54), .S(sum[9]) );
  ADDHXL U59 ( .A(a[7]), .B(n57), .CO(n56), .S(sum[7]) );
  ADDHXL U62 ( .A(a[4]), .B(n60), .CO(n59), .S(sum[4]) );
  ADDHXL U64 ( .A(a[2]), .B(n62), .CO(n61), .S(sum[2]) );
  ADDHXL U66 ( .A(carry_in), .B(a[0]), .CO(n63), .S(sum[0]) );
  ADDHXL U70 ( .A(a[47]), .B(n17), .CO(n16), .S(sum[47]) );
  ADDHXL U71 ( .A(a[44]), .B(n20), .CO(n19), .S(sum[44]) );
  ADDHXL U72 ( .A(a[55]), .B(n9), .CO(n8), .S(sum[55]) );
  ADDHXL U73 ( .A(a[46]), .B(n18), .CO(n17), .S(sum[46]) );
  ADDHXL U74 ( .A(a[43]), .B(n21), .CO(n20), .S(sum[43]) );
  ADDHXL U75 ( .A(a[54]), .B(n10), .CO(n9), .S(sum[54]) );
  ADDHX2 U76 ( .A(a[59]), .B(n5), .CO(n4), .S(sum[59]) );
  ADDHX1 U77 ( .A(a[38]), .B(n26), .CO(n25), .S(sum[38]) );
  ADDHX1 U78 ( .A(a[33]), .B(n31), .CO(n30), .S(sum[33]) );
  ADDHX1 U79 ( .A(a[22]), .B(n42), .CO(n41), .S(sum[22]) );
  ADDHX1 U80 ( .A(a[20]), .B(n44), .CO(n43), .S(sum[20]) );
  ADDHX1 U81 ( .A(a[51]), .B(n13), .CO(n12), .S(sum[51]) );
  ADDHX1 U82 ( .A(a[49]), .B(n15), .CO(n14), .S(sum[49]) );
  ADDHX1 U83 ( .A(a[40]), .B(n24), .CO(n23), .S(sum[40]) );
  ADDHX1 U84 ( .A(a[35]), .B(n29), .CO(n28), .S(sum[35]) );
  ADDHX1 U85 ( .A(a[28]), .B(n36), .CO(n35), .S(sum[28]) );
  ADDHX1 U86 ( .A(a[25]), .B(n39), .CO(n38), .S(sum[25]) );
  ADDHX1 U87 ( .A(a[15]), .B(n49), .CO(n48), .S(sum[15]) );
  ADDHX1 U88 ( .A(a[10]), .B(n54), .CO(n53), .S(sum[10]) );
  ADDHX1 U89 ( .A(a[3]), .B(n61), .CO(n60), .S(sum[3]) );
  ADDHX1 U90 ( .A(a[8]), .B(n56), .CO(n55), .S(sum[8]) );
  ADDHX1 U91 ( .A(a[1]), .B(n63), .CO(n62), .S(sum[1]) );
  ADDHX1 U92 ( .A(a[57]), .B(n7), .CO(n6), .S(sum[57]) );
  ADDHX1 U93 ( .A(a[31]), .B(n33), .CO(n32), .S(sum[31]) );
  ADDHX1 U94 ( .A(a[13]), .B(n51), .CO(n50), .S(sum[13]) );
  ADDHX1 U95 ( .A(a[5]), .B(n59), .CO(n58), .S(sum[5]) );
  ADDHX1 U96 ( .A(a[18]), .B(n46), .CO(n45), .S(sum[18]) );
  ADDHXL U97 ( .A(a[52]), .B(n12), .CO(n11), .S(sum[52]) );
  ADDHXL U98 ( .A(a[41]), .B(n23), .CO(n22), .S(sum[41]) );
  ADDHXL U99 ( .A(a[16]), .B(n48), .CO(n47), .S(sum[16]) );
  ADDHXL U100 ( .A(a[23]), .B(n41), .CO(n40), .S(sum[23]) );
  ADDHXL U101 ( .A(a[26]), .B(n38), .CO(n37), .S(sum[26]) );
  ADDHXL U102 ( .A(a[36]), .B(n28), .CO(n27), .S(sum[36]) );
  ADDHXL U103 ( .A(a[29]), .B(n35), .CO(n34), .S(sum[29]) );
  XOR2XL U104 ( .A(n4), .B(a[60]), .Y(sum[60]) );
  ADDHXL U105 ( .A(a[17]), .B(n47), .CO(n46), .S(sum[17]) );
  ADDHXL U106 ( .A(a[6]), .B(n58), .CO(n57), .S(sum[6]) );
  ADDHXL U107 ( .A(a[14]), .B(n50), .CO(n49), .S(sum[14]) );
  ADDHXL U108 ( .A(a[32]), .B(n32), .CO(n31), .S(sum[32]) );
  NOR2BX1 U109 ( .AN(a[60]), .B(n4), .Y(\sum[63] ) );
endmodule


module GSIM_DW_div_tc_2 ( a, b, quotient, remainder, divide_by_0 );
  input [63:0] a;
  input [5:0] b;
  output [63:0] quotient;
  output [5:0] remainder;
  output divide_by_0;
  wire   \u_div/QInv[63] , \u_div/QInv[59] , \u_div/QInv[58] ,
         \u_div/QInv[57] , \u_div/QInv[56] , \u_div/QInv[55] ,
         \u_div/QInv[54] , \u_div/QInv[53] , \u_div/QInv[52] ,
         \u_div/QInv[51] , \u_div/QInv[50] , \u_div/QInv[49] ,
         \u_div/QInv[48] , \u_div/QInv[47] , \u_div/QInv[46] ,
         \u_div/QInv[45] , \u_div/QInv[44] , \u_div/QInv[43] ,
         \u_div/QInv[42] , \u_div/QInv[41] , \u_div/QInv[40] ,
         \u_div/QInv[39] , \u_div/QInv[38] , \u_div/QInv[37] ,
         \u_div/QInv[36] , \u_div/QInv[35] , \u_div/QInv[34] ,
         \u_div/QInv[33] , \u_div/QInv[32] , \u_div/QInv[31] ,
         \u_div/QInv[30] , \u_div/QInv[29] , \u_div/QInv[28] ,
         \u_div/QInv[27] , \u_div/QInv[26] , \u_div/QInv[25] ,
         \u_div/QInv[24] , \u_div/QInv[23] , \u_div/QInv[22] ,
         \u_div/QInv[21] , \u_div/QInv[20] , \u_div/QInv[19] ,
         \u_div/QInv[18] , \u_div/QInv[17] , \u_div/QInv[16] ,
         \u_div/QInv[15] , \u_div/QInv[14] , \u_div/QInv[13] ,
         \u_div/QInv[12] , \u_div/QInv[11] , \u_div/QInv[10] , \u_div/QInv[9] ,
         \u_div/QInv[8] , \u_div/QInv[7] , \u_div/QInv[6] , \u_div/QInv[5] ,
         \u_div/QInv[4] , \u_div/QInv[3] , \u_div/QInv[2] , \u_div/QInv[1] ,
         \u_div/QInv[0] , \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] ,
         \u_div/SumTmp[1][3] , \u_div/SumTmp[1][4] , \u_div/SumTmp[2][1] ,
         \u_div/SumTmp[2][2] , \u_div/SumTmp[2][3] , \u_div/SumTmp[2][4] ,
         \u_div/SumTmp[3][1] , \u_div/SumTmp[3][2] , \u_div/SumTmp[3][3] ,
         \u_div/SumTmp[3][4] , \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] ,
         \u_div/SumTmp[4][3] , \u_div/SumTmp[4][4] , \u_div/SumTmp[5][1] ,
         \u_div/SumTmp[5][2] , \u_div/SumTmp[5][3] , \u_div/SumTmp[5][4] ,
         \u_div/SumTmp[6][1] , \u_div/SumTmp[6][2] , \u_div/SumTmp[6][3] ,
         \u_div/SumTmp[6][4] , \u_div/SumTmp[7][1] , \u_div/SumTmp[7][2] ,
         \u_div/SumTmp[7][3] , \u_div/SumTmp[7][4] , \u_div/SumTmp[8][1] ,
         \u_div/SumTmp[8][2] , \u_div/SumTmp[8][3] , \u_div/SumTmp[8][4] ,
         \u_div/SumTmp[9][1] , \u_div/SumTmp[9][2] , \u_div/SumTmp[9][3] ,
         \u_div/SumTmp[9][4] , \u_div/SumTmp[10][1] , \u_div/SumTmp[10][2] ,
         \u_div/SumTmp[10][3] , \u_div/SumTmp[10][4] , \u_div/SumTmp[11][1] ,
         \u_div/SumTmp[11][2] , \u_div/SumTmp[11][3] , \u_div/SumTmp[11][4] ,
         \u_div/SumTmp[12][1] , \u_div/SumTmp[12][2] , \u_div/SumTmp[12][3] ,
         \u_div/SumTmp[12][4] , \u_div/SumTmp[13][1] , \u_div/SumTmp[13][2] ,
         \u_div/SumTmp[13][3] , \u_div/SumTmp[13][4] , \u_div/SumTmp[14][1] ,
         \u_div/SumTmp[14][2] , \u_div/SumTmp[14][3] , \u_div/SumTmp[14][4] ,
         \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] , \u_div/SumTmp[15][3] ,
         \u_div/SumTmp[15][4] , \u_div/SumTmp[16][1] , \u_div/SumTmp[16][2] ,
         \u_div/SumTmp[16][3] , \u_div/SumTmp[16][4] , \u_div/SumTmp[17][1] ,
         \u_div/SumTmp[17][2] , \u_div/SumTmp[17][3] , \u_div/SumTmp[17][4] ,
         \u_div/SumTmp[18][1] , \u_div/SumTmp[18][2] , \u_div/SumTmp[18][3] ,
         \u_div/SumTmp[18][4] , \u_div/SumTmp[19][1] , \u_div/SumTmp[19][2] ,
         \u_div/SumTmp[19][3] , \u_div/SumTmp[19][4] , \u_div/SumTmp[20][1] ,
         \u_div/SumTmp[20][2] , \u_div/SumTmp[20][3] , \u_div/SumTmp[20][4] ,
         \u_div/SumTmp[21][1] , \u_div/SumTmp[21][2] , \u_div/SumTmp[21][3] ,
         \u_div/SumTmp[21][4] , \u_div/SumTmp[22][1] , \u_div/SumTmp[22][2] ,
         \u_div/SumTmp[22][3] , \u_div/SumTmp[22][4] , \u_div/SumTmp[23][1] ,
         \u_div/SumTmp[23][2] , \u_div/SumTmp[23][3] , \u_div/SumTmp[23][4] ,
         \u_div/SumTmp[24][1] , \u_div/SumTmp[24][2] , \u_div/SumTmp[24][3] ,
         \u_div/SumTmp[24][4] , \u_div/SumTmp[25][1] , \u_div/SumTmp[25][2] ,
         \u_div/SumTmp[25][3] , \u_div/SumTmp[25][4] , \u_div/SumTmp[26][1] ,
         \u_div/SumTmp[26][2] , \u_div/SumTmp[26][3] , \u_div/SumTmp[26][4] ,
         \u_div/SumTmp[27][1] , \u_div/SumTmp[27][2] , \u_div/SumTmp[27][3] ,
         \u_div/SumTmp[27][4] , \u_div/SumTmp[28][1] , \u_div/SumTmp[28][2] ,
         \u_div/SumTmp[28][3] , \u_div/SumTmp[28][4] , \u_div/SumTmp[29][1] ,
         \u_div/SumTmp[29][2] , \u_div/SumTmp[29][3] , \u_div/SumTmp[29][4] ,
         \u_div/SumTmp[30][1] , \u_div/SumTmp[30][2] , \u_div/SumTmp[30][3] ,
         \u_div/SumTmp[30][4] , \u_div/SumTmp[31][1] , \u_div/SumTmp[31][2] ,
         \u_div/SumTmp[31][3] , \u_div/SumTmp[31][4] , \u_div/SumTmp[32][1] ,
         \u_div/SumTmp[32][2] , \u_div/SumTmp[32][3] , \u_div/SumTmp[32][4] ,
         \u_div/SumTmp[33][1] , \u_div/SumTmp[33][2] , \u_div/SumTmp[33][3] ,
         \u_div/SumTmp[33][4] , \u_div/SumTmp[34][1] , \u_div/SumTmp[34][2] ,
         \u_div/SumTmp[34][3] , \u_div/SumTmp[34][4] , \u_div/SumTmp[35][1] ,
         \u_div/SumTmp[35][2] , \u_div/SumTmp[35][3] , \u_div/SumTmp[35][4] ,
         \u_div/SumTmp[36][1] , \u_div/SumTmp[36][2] , \u_div/SumTmp[36][3] ,
         \u_div/SumTmp[36][4] , \u_div/SumTmp[37][1] , \u_div/SumTmp[37][2] ,
         \u_div/SumTmp[37][3] , \u_div/SumTmp[37][4] , \u_div/SumTmp[38][1] ,
         \u_div/SumTmp[38][2] , \u_div/SumTmp[38][3] , \u_div/SumTmp[38][4] ,
         \u_div/SumTmp[39][1] , \u_div/SumTmp[39][2] , \u_div/SumTmp[39][3] ,
         \u_div/SumTmp[39][4] , \u_div/SumTmp[40][1] , \u_div/SumTmp[40][2] ,
         \u_div/SumTmp[40][3] , \u_div/SumTmp[40][4] , \u_div/SumTmp[41][1] ,
         \u_div/SumTmp[41][2] , \u_div/SumTmp[41][3] , \u_div/SumTmp[41][4] ,
         \u_div/SumTmp[42][1] , \u_div/SumTmp[42][2] , \u_div/SumTmp[42][3] ,
         \u_div/SumTmp[42][4] , \u_div/SumTmp[43][1] , \u_div/SumTmp[43][2] ,
         \u_div/SumTmp[43][3] , \u_div/SumTmp[43][4] , \u_div/SumTmp[44][1] ,
         \u_div/SumTmp[44][2] , \u_div/SumTmp[44][3] , \u_div/SumTmp[44][4] ,
         \u_div/SumTmp[45][1] , \u_div/SumTmp[45][2] , \u_div/SumTmp[45][3] ,
         \u_div/SumTmp[45][4] , \u_div/SumTmp[46][1] , \u_div/SumTmp[46][2] ,
         \u_div/SumTmp[46][3] , \u_div/SumTmp[46][4] , \u_div/SumTmp[47][1] ,
         \u_div/SumTmp[47][2] , \u_div/SumTmp[47][3] , \u_div/SumTmp[47][4] ,
         \u_div/SumTmp[48][1] , \u_div/SumTmp[48][2] , \u_div/SumTmp[48][3] ,
         \u_div/SumTmp[48][4] , \u_div/SumTmp[49][1] , \u_div/SumTmp[49][2] ,
         \u_div/SumTmp[49][3] , \u_div/SumTmp[49][4] , \u_div/SumTmp[50][1] ,
         \u_div/SumTmp[50][2] , \u_div/SumTmp[50][3] , \u_div/SumTmp[50][4] ,
         \u_div/SumTmp[51][1] , \u_div/SumTmp[51][2] , \u_div/SumTmp[51][3] ,
         \u_div/SumTmp[51][4] , \u_div/SumTmp[52][1] , \u_div/SumTmp[52][2] ,
         \u_div/SumTmp[52][3] , \u_div/SumTmp[52][4] , \u_div/SumTmp[53][1] ,
         \u_div/SumTmp[53][2] , \u_div/SumTmp[53][3] , \u_div/SumTmp[53][4] ,
         \u_div/SumTmp[54][1] , \u_div/SumTmp[54][2] , \u_div/SumTmp[54][3] ,
         \u_div/SumTmp[54][4] , \u_div/SumTmp[55][1] , \u_div/SumTmp[55][2] ,
         \u_div/SumTmp[55][3] , \u_div/SumTmp[55][4] , \u_div/SumTmp[56][1] ,
         \u_div/SumTmp[56][2] , \u_div/SumTmp[56][3] , \u_div/SumTmp[56][4] ,
         \u_div/SumTmp[57][1] , \u_div/SumTmp[57][2] , \u_div/SumTmp[57][3] ,
         \u_div/SumTmp[57][4] , \u_div/SumTmp[58][1] , \u_div/SumTmp[58][2] ,
         \u_div/SumTmp[58][3] , \u_div/SumTmp[58][4] , \u_div/SumTmp[59][3] ,
         \u_div/SumTmp[59][4] , \u_div/CryTmp[0][6] , \u_div/CryTmp[1][6] ,
         \u_div/CryTmp[2][6] , \u_div/CryTmp[3][6] , \u_div/CryTmp[4][6] ,
         \u_div/CryTmp[5][6] , \u_div/CryTmp[6][6] , \u_div/CryTmp[7][6] ,
         \u_div/CryTmp[8][6] , \u_div/CryTmp[9][6] , \u_div/CryTmp[10][6] ,
         \u_div/CryTmp[11][6] , \u_div/CryTmp[12][6] , \u_div/CryTmp[13][6] ,
         \u_div/CryTmp[14][6] , \u_div/CryTmp[15][6] , \u_div/CryTmp[16][6] ,
         \u_div/CryTmp[17][6] , \u_div/CryTmp[18][6] , \u_div/CryTmp[19][6] ,
         \u_div/CryTmp[20][6] , \u_div/CryTmp[21][6] , \u_div/CryTmp[22][6] ,
         \u_div/CryTmp[23][6] , \u_div/CryTmp[24][6] , \u_div/CryTmp[25][6] ,
         \u_div/CryTmp[26][6] , \u_div/CryTmp[27][6] , \u_div/CryTmp[28][6] ,
         \u_div/CryTmp[29][6] , \u_div/CryTmp[30][6] , \u_div/CryTmp[31][6] ,
         \u_div/CryTmp[32][6] , \u_div/CryTmp[33][6] , \u_div/CryTmp[34][6] ,
         \u_div/CryTmp[35][6] , \u_div/CryTmp[36][6] , \u_div/CryTmp[37][6] ,
         \u_div/CryTmp[38][6] , \u_div/CryTmp[39][6] , \u_div/CryTmp[40][6] ,
         \u_div/CryTmp[41][6] , \u_div/CryTmp[42][6] , \u_div/CryTmp[43][6] ,
         \u_div/CryTmp[44][6] , \u_div/CryTmp[45][6] , \u_div/CryTmp[46][6] ,
         \u_div/CryTmp[47][6] , \u_div/CryTmp[48][6] , \u_div/CryTmp[49][6] ,
         \u_div/CryTmp[50][6] , \u_div/CryTmp[51][6] , \u_div/CryTmp[52][6] ,
         \u_div/CryTmp[53][6] , \u_div/CryTmp[54][6] , \u_div/CryTmp[55][6] ,
         \u_div/CryTmp[56][6] , \u_div/CryTmp[57][6] , \u_div/CryTmp[58][6] ,
         \u_div/CryTmp[59][6] , \u_div/PartRem[1][3] , \u_div/PartRem[1][4] ,
         \u_div/PartRem[1][5] , \u_div/PartRem[2][2] , \u_div/PartRem[2][3] ,
         \u_div/PartRem[2][4] , \u_div/PartRem[2][5] , \u_div/PartRem[3][0] ,
         \u_div/PartRem[3][2] , \u_div/PartRem[3][3] , \u_div/PartRem[3][4] ,
         \u_div/PartRem[3][5] , \u_div/PartRem[4][0] , \u_div/PartRem[4][2] ,
         \u_div/PartRem[4][3] , \u_div/PartRem[4][4] , \u_div/PartRem[4][5] ,
         \u_div/PartRem[5][0] , \u_div/PartRem[5][2] , \u_div/PartRem[5][3] ,
         \u_div/PartRem[5][4] , \u_div/PartRem[5][5] , \u_div/PartRem[6][0] ,
         \u_div/PartRem[6][2] , \u_div/PartRem[6][3] , \u_div/PartRem[6][4] ,
         \u_div/PartRem[6][5] , \u_div/PartRem[7][0] , \u_div/PartRem[7][2] ,
         \u_div/PartRem[7][3] , \u_div/PartRem[7][4] , \u_div/PartRem[7][5] ,
         \u_div/PartRem[8][0] , \u_div/PartRem[8][2] , \u_div/PartRem[8][3] ,
         \u_div/PartRem[8][4] , \u_div/PartRem[8][5] , \u_div/PartRem[9][0] ,
         \u_div/PartRem[9][2] , \u_div/PartRem[9][3] , \u_div/PartRem[9][4] ,
         \u_div/PartRem[9][5] , \u_div/PartRem[10][0] , \u_div/PartRem[10][2] ,
         \u_div/PartRem[10][3] , \u_div/PartRem[10][4] ,
         \u_div/PartRem[10][5] , \u_div/PartRem[11][0] ,
         \u_div/PartRem[11][2] , \u_div/PartRem[11][3] ,
         \u_div/PartRem[11][4] , \u_div/PartRem[11][5] ,
         \u_div/PartRem[12][0] , \u_div/PartRem[12][2] ,
         \u_div/PartRem[12][3] , \u_div/PartRem[12][4] ,
         \u_div/PartRem[12][5] , \u_div/PartRem[13][0] ,
         \u_div/PartRem[13][2] , \u_div/PartRem[13][3] ,
         \u_div/PartRem[13][4] , \u_div/PartRem[13][5] ,
         \u_div/PartRem[14][0] , \u_div/PartRem[14][2] ,
         \u_div/PartRem[14][3] , \u_div/PartRem[14][4] ,
         \u_div/PartRem[14][5] , \u_div/PartRem[15][0] ,
         \u_div/PartRem[15][2] , \u_div/PartRem[15][3] ,
         \u_div/PartRem[15][4] , \u_div/PartRem[15][5] ,
         \u_div/PartRem[16][0] , \u_div/PartRem[16][2] ,
         \u_div/PartRem[16][3] , \u_div/PartRem[16][4] ,
         \u_div/PartRem[16][5] , \u_div/PartRem[17][0] ,
         \u_div/PartRem[17][2] , \u_div/PartRem[17][3] ,
         \u_div/PartRem[17][4] , \u_div/PartRem[17][5] ,
         \u_div/PartRem[18][0] , \u_div/PartRem[18][2] ,
         \u_div/PartRem[18][3] , \u_div/PartRem[18][4] ,
         \u_div/PartRem[18][5] , \u_div/PartRem[19][0] ,
         \u_div/PartRem[19][2] , \u_div/PartRem[19][3] ,
         \u_div/PartRem[19][4] , \u_div/PartRem[19][5] ,
         \u_div/PartRem[20][0] , \u_div/PartRem[20][2] ,
         \u_div/PartRem[20][3] , \u_div/PartRem[20][4] ,
         \u_div/PartRem[20][5] , \u_div/PartRem[21][0] ,
         \u_div/PartRem[21][2] , \u_div/PartRem[21][3] ,
         \u_div/PartRem[21][4] , \u_div/PartRem[21][5] ,
         \u_div/PartRem[22][0] , \u_div/PartRem[22][2] ,
         \u_div/PartRem[22][3] , \u_div/PartRem[22][4] ,
         \u_div/PartRem[22][5] , \u_div/PartRem[23][0] ,
         \u_div/PartRem[23][2] , \u_div/PartRem[23][3] ,
         \u_div/PartRem[23][4] , \u_div/PartRem[23][5] ,
         \u_div/PartRem[24][0] , \u_div/PartRem[24][2] ,
         \u_div/PartRem[24][3] , \u_div/PartRem[24][4] ,
         \u_div/PartRem[24][5] , \u_div/PartRem[25][0] ,
         \u_div/PartRem[25][2] , \u_div/PartRem[25][3] ,
         \u_div/PartRem[25][4] , \u_div/PartRem[25][5] ,
         \u_div/PartRem[26][0] , \u_div/PartRem[26][2] ,
         \u_div/PartRem[26][3] , \u_div/PartRem[26][4] ,
         \u_div/PartRem[26][5] , \u_div/PartRem[27][0] ,
         \u_div/PartRem[27][2] , \u_div/PartRem[27][3] ,
         \u_div/PartRem[27][4] , \u_div/PartRem[27][5] ,
         \u_div/PartRem[28][0] , \u_div/PartRem[28][2] ,
         \u_div/PartRem[28][3] , \u_div/PartRem[28][4] ,
         \u_div/PartRem[28][5] , \u_div/PartRem[29][0] ,
         \u_div/PartRem[29][2] , \u_div/PartRem[29][3] ,
         \u_div/PartRem[29][4] , \u_div/PartRem[29][5] ,
         \u_div/PartRem[30][0] , \u_div/PartRem[30][2] ,
         \u_div/PartRem[30][3] , \u_div/PartRem[30][4] ,
         \u_div/PartRem[30][5] , \u_div/PartRem[31][0] ,
         \u_div/PartRem[31][2] , \u_div/PartRem[31][3] ,
         \u_div/PartRem[31][4] , \u_div/PartRem[31][5] ,
         \u_div/PartRem[32][0] , \u_div/PartRem[32][2] ,
         \u_div/PartRem[32][3] , \u_div/PartRem[32][4] ,
         \u_div/PartRem[32][5] , \u_div/PartRem[33][0] ,
         \u_div/PartRem[33][2] , \u_div/PartRem[33][3] ,
         \u_div/PartRem[33][4] , \u_div/PartRem[33][5] ,
         \u_div/PartRem[34][0] , \u_div/PartRem[34][2] ,
         \u_div/PartRem[34][3] , \u_div/PartRem[34][4] ,
         \u_div/PartRem[34][5] , \u_div/PartRem[35][0] ,
         \u_div/PartRem[35][2] , \u_div/PartRem[35][3] ,
         \u_div/PartRem[35][4] , \u_div/PartRem[35][5] ,
         \u_div/PartRem[36][0] , \u_div/PartRem[36][2] ,
         \u_div/PartRem[36][3] , \u_div/PartRem[36][4] ,
         \u_div/PartRem[36][5] , \u_div/PartRem[37][0] ,
         \u_div/PartRem[37][2] , \u_div/PartRem[37][3] ,
         \u_div/PartRem[37][4] , \u_div/PartRem[37][5] ,
         \u_div/PartRem[38][0] , \u_div/PartRem[38][2] ,
         \u_div/PartRem[38][3] , \u_div/PartRem[38][4] ,
         \u_div/PartRem[38][5] , \u_div/PartRem[39][0] ,
         \u_div/PartRem[39][2] , \u_div/PartRem[39][3] ,
         \u_div/PartRem[39][4] , \u_div/PartRem[39][5] ,
         \u_div/PartRem[40][0] , \u_div/PartRem[40][2] ,
         \u_div/PartRem[40][3] , \u_div/PartRem[40][4] ,
         \u_div/PartRem[40][5] , \u_div/PartRem[41][0] ,
         \u_div/PartRem[41][2] , \u_div/PartRem[41][3] ,
         \u_div/PartRem[41][4] , \u_div/PartRem[41][5] ,
         \u_div/PartRem[42][0] , \u_div/PartRem[42][2] ,
         \u_div/PartRem[42][3] , \u_div/PartRem[42][4] ,
         \u_div/PartRem[42][5] , \u_div/PartRem[43][0] ,
         \u_div/PartRem[43][2] , \u_div/PartRem[43][3] ,
         \u_div/PartRem[43][4] , \u_div/PartRem[43][5] ,
         \u_div/PartRem[44][0] , \u_div/PartRem[44][2] ,
         \u_div/PartRem[44][3] , \u_div/PartRem[44][4] ,
         \u_div/PartRem[44][5] , \u_div/PartRem[45][0] ,
         \u_div/PartRem[45][2] , \u_div/PartRem[45][3] ,
         \u_div/PartRem[45][4] , \u_div/PartRem[45][5] ,
         \u_div/PartRem[46][0] , \u_div/PartRem[46][2] ,
         \u_div/PartRem[46][3] , \u_div/PartRem[46][4] ,
         \u_div/PartRem[46][5] , \u_div/PartRem[47][0] ,
         \u_div/PartRem[47][2] , \u_div/PartRem[47][3] ,
         \u_div/PartRem[47][4] , \u_div/PartRem[47][5] ,
         \u_div/PartRem[48][0] , \u_div/PartRem[48][2] ,
         \u_div/PartRem[48][3] , \u_div/PartRem[48][4] ,
         \u_div/PartRem[48][5] , \u_div/PartRem[49][0] ,
         \u_div/PartRem[49][2] , \u_div/PartRem[49][3] ,
         \u_div/PartRem[49][4] , \u_div/PartRem[49][5] ,
         \u_div/PartRem[50][0] , \u_div/PartRem[50][2] ,
         \u_div/PartRem[50][3] , \u_div/PartRem[50][4] ,
         \u_div/PartRem[50][5] , \u_div/PartRem[51][0] ,
         \u_div/PartRem[51][2] , \u_div/PartRem[51][3] ,
         \u_div/PartRem[51][4] , \u_div/PartRem[51][5] ,
         \u_div/PartRem[52][0] , \u_div/PartRem[52][2] ,
         \u_div/PartRem[52][3] , \u_div/PartRem[52][4] ,
         \u_div/PartRem[52][5] , \u_div/PartRem[53][0] ,
         \u_div/PartRem[53][2] , \u_div/PartRem[53][3] ,
         \u_div/PartRem[53][4] , \u_div/PartRem[53][5] ,
         \u_div/PartRem[54][0] , \u_div/PartRem[54][2] ,
         \u_div/PartRem[54][3] , \u_div/PartRem[54][4] ,
         \u_div/PartRem[54][5] , \u_div/PartRem[55][0] ,
         \u_div/PartRem[55][2] , \u_div/PartRem[55][3] ,
         \u_div/PartRem[55][4] , \u_div/PartRem[55][5] ,
         \u_div/PartRem[56][0] , \u_div/PartRem[56][2] ,
         \u_div/PartRem[56][3] , \u_div/PartRem[56][4] ,
         \u_div/PartRem[56][5] , \u_div/PartRem[57][0] ,
         \u_div/PartRem[57][2] , \u_div/PartRem[57][3] ,
         \u_div/PartRem[57][4] , \u_div/PartRem[57][5] ,
         \u_div/PartRem[58][0] , \u_div/PartRem[58][2] ,
         \u_div/PartRem[58][3] , \u_div/PartRem[58][4] ,
         \u_div/PartRem[58][5] , \u_div/PartRem[59][0] ,
         \u_div/PartRem[59][2] , \u_div/PartRem[59][3] ,
         \u_div/PartRem[59][4] , \u_div/PartRem[59][5] ,
         \u_div/PartRem[60][0] , \u_div/PartRem[61][0] ,
         \u_div/PartRem[62][0] , \u_div/PartRem[63][0] ,
         \u_div/PartRem[64][0] , \u_div/u_add_PartRem_2_1/n3 ,
         \u_div/u_add_PartRem_2_1/n2 , \u_div/u_add_PartRem_2_2/n3 ,
         \u_div/u_add_PartRem_2_2/n2 , \u_div/u_add_PartRem_2_3/n3 ,
         \u_div/u_add_PartRem_2_3/n2 , \u_div/u_add_PartRem_2_4/n3 ,
         \u_div/u_add_PartRem_2_4/n2 , \u_div/u_add_PartRem_2_5/n3 ,
         \u_div/u_add_PartRem_2_5/n2 , \u_div/u_add_PartRem_2_6/n3 ,
         \u_div/u_add_PartRem_2_6/n2 , \u_div/u_add_PartRem_2_7/n3 ,
         \u_div/u_add_PartRem_2_7/n2 , \u_div/u_add_PartRem_2_8/n3 ,
         \u_div/u_add_PartRem_2_8/n2 , \u_div/u_add_PartRem_2_9/n3 ,
         \u_div/u_add_PartRem_2_9/n2 , \u_div/u_add_PartRem_2_10/n3 ,
         \u_div/u_add_PartRem_2_10/n2 , \u_div/u_add_PartRem_2_11/n3 ,
         \u_div/u_add_PartRem_2_11/n2 , \u_div/u_add_PartRem_2_12/n3 ,
         \u_div/u_add_PartRem_2_12/n2 , \u_div/u_add_PartRem_2_13/n3 ,
         \u_div/u_add_PartRem_2_13/n2 , \u_div/u_add_PartRem_2_14/n3 ,
         \u_div/u_add_PartRem_2_14/n2 , \u_div/u_add_PartRem_2_15/n3 ,
         \u_div/u_add_PartRem_2_15/n2 , \u_div/u_add_PartRem_2_16/n3 ,
         \u_div/u_add_PartRem_2_16/n2 , \u_div/u_add_PartRem_2_17/n3 ,
         \u_div/u_add_PartRem_2_17/n2 , \u_div/u_add_PartRem_2_18/n3 ,
         \u_div/u_add_PartRem_2_18/n2 , \u_div/u_add_PartRem_2_19/n3 ,
         \u_div/u_add_PartRem_2_19/n2 , \u_div/u_add_PartRem_2_20/n3 ,
         \u_div/u_add_PartRem_2_20/n2 , \u_div/u_add_PartRem_2_21/n3 ,
         \u_div/u_add_PartRem_2_21/n2 , \u_div/u_add_PartRem_2_22/n3 ,
         \u_div/u_add_PartRem_2_22/n2 , \u_div/u_add_PartRem_2_23/n3 ,
         \u_div/u_add_PartRem_2_23/n2 , \u_div/u_add_PartRem_2_24/n3 ,
         \u_div/u_add_PartRem_2_24/n2 , \u_div/u_add_PartRem_2_25/n3 ,
         \u_div/u_add_PartRem_2_25/n2 , \u_div/u_add_PartRem_2_26/n3 ,
         \u_div/u_add_PartRem_2_26/n2 , \u_div/u_add_PartRem_2_27/n3 ,
         \u_div/u_add_PartRem_2_27/n2 , \u_div/u_add_PartRem_2_28/n3 ,
         \u_div/u_add_PartRem_2_28/n2 , \u_div/u_add_PartRem_2_29/n3 ,
         \u_div/u_add_PartRem_2_29/n2 , \u_div/u_add_PartRem_2_30/n3 ,
         \u_div/u_add_PartRem_2_30/n2 , \u_div/u_add_PartRem_2_31/n3 ,
         \u_div/u_add_PartRem_2_31/n2 , \u_div/u_add_PartRem_2_32/n3 ,
         \u_div/u_add_PartRem_2_32/n2 , \u_div/u_add_PartRem_2_33/n3 ,
         \u_div/u_add_PartRem_2_33/n2 , \u_div/u_add_PartRem_2_34/n3 ,
         \u_div/u_add_PartRem_2_34/n2 , \u_div/u_add_PartRem_2_35/n3 ,
         \u_div/u_add_PartRem_2_35/n2 , \u_div/u_add_PartRem_2_36/n3 ,
         \u_div/u_add_PartRem_2_36/n2 , \u_div/u_add_PartRem_2_37/n3 ,
         \u_div/u_add_PartRem_2_37/n2 , \u_div/u_add_PartRem_2_38/n3 ,
         \u_div/u_add_PartRem_2_38/n2 , \u_div/u_add_PartRem_2_39/n3 ,
         \u_div/u_add_PartRem_2_39/n2 , \u_div/u_add_PartRem_2_40/n3 ,
         \u_div/u_add_PartRem_2_40/n2 , \u_div/u_add_PartRem_2_41/n3 ,
         \u_div/u_add_PartRem_2_41/n2 , \u_div/u_add_PartRem_2_42/n3 ,
         \u_div/u_add_PartRem_2_42/n2 , \u_div/u_add_PartRem_2_43/n3 ,
         \u_div/u_add_PartRem_2_43/n2 , \u_div/u_add_PartRem_2_44/n3 ,
         \u_div/u_add_PartRem_2_44/n2 , \u_div/u_add_PartRem_2_45/n3 ,
         \u_div/u_add_PartRem_2_45/n2 , \u_div/u_add_PartRem_2_46/n3 ,
         \u_div/u_add_PartRem_2_46/n2 , \u_div/u_add_PartRem_2_47/n3 ,
         \u_div/u_add_PartRem_2_47/n2 , \u_div/u_add_PartRem_2_48/n3 ,
         \u_div/u_add_PartRem_2_48/n2 , \u_div/u_add_PartRem_2_49/n3 ,
         \u_div/u_add_PartRem_2_49/n2 , \u_div/u_add_PartRem_2_50/n3 ,
         \u_div/u_add_PartRem_2_50/n2 , \u_div/u_add_PartRem_2_51/n3 ,
         \u_div/u_add_PartRem_2_51/n2 , \u_div/u_add_PartRem_2_52/n3 ,
         \u_div/u_add_PartRem_2_52/n2 , \u_div/u_add_PartRem_2_53/n3 ,
         \u_div/u_add_PartRem_2_53/n2 , \u_div/u_add_PartRem_2_54/n3 ,
         \u_div/u_add_PartRem_2_54/n2 , \u_div/u_add_PartRem_2_55/n3 ,
         \u_div/u_add_PartRem_2_55/n2 , \u_div/u_add_PartRem_2_56/n3 ,
         \u_div/u_add_PartRem_2_56/n2 , \u_div/u_add_PartRem_2_57/n3 ,
         \u_div/u_add_PartRem_2_57/n2 , \u_div/u_add_PartRem_2_58/n3 ,
         \u_div/u_add_PartRem_2_58/n2 , n1, n2, n3, n4, n5, n6, n7, n8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign \u_div/QInv[63]  = a[63];

  GSIM_DW01_absval_2 \u_div/u_absval_AAbs  ( .A({n3, a[62:0]}), .ABSVAL({
        \u_div/PartRem[64][0] , \u_div/PartRem[63][0] , \u_div/PartRem[62][0] , 
        \u_div/PartRem[61][0] , \u_div/PartRem[60][0] , \u_div/PartRem[59][0] , 
        \u_div/PartRem[58][0] , \u_div/PartRem[57][0] , \u_div/PartRem[56][0] , 
        \u_div/PartRem[55][0] , \u_div/PartRem[54][0] , \u_div/PartRem[53][0] , 
        \u_div/PartRem[52][0] , \u_div/PartRem[51][0] , \u_div/PartRem[50][0] , 
        \u_div/PartRem[49][0] , \u_div/PartRem[48][0] , \u_div/PartRem[47][0] , 
        \u_div/PartRem[46][0] , \u_div/PartRem[45][0] , \u_div/PartRem[44][0] , 
        \u_div/PartRem[43][0] , \u_div/PartRem[42][0] , \u_div/PartRem[41][0] , 
        \u_div/PartRem[40][0] , \u_div/PartRem[39][0] , \u_div/PartRem[38][0] , 
        \u_div/PartRem[37][0] , \u_div/PartRem[36][0] , \u_div/PartRem[35][0] , 
        \u_div/PartRem[34][0] , \u_div/PartRem[33][0] , \u_div/PartRem[32][0] , 
        \u_div/PartRem[31][0] , \u_div/PartRem[30][0] , \u_div/PartRem[29][0] , 
        \u_div/PartRem[28][0] , \u_div/PartRem[27][0] , \u_div/PartRem[26][0] , 
        \u_div/PartRem[25][0] , \u_div/PartRem[24][0] , \u_div/PartRem[23][0] , 
        \u_div/PartRem[22][0] , \u_div/PartRem[21][0] , \u_div/PartRem[20][0] , 
        \u_div/PartRem[19][0] , \u_div/PartRem[18][0] , \u_div/PartRem[17][0] , 
        \u_div/PartRem[16][0] , \u_div/PartRem[15][0] , \u_div/PartRem[14][0] , 
        \u_div/PartRem[13][0] , \u_div/PartRem[12][0] , \u_div/PartRem[11][0] , 
        \u_div/PartRem[10][0] , \u_div/PartRem[9][0] , \u_div/PartRem[8][0] , 
        \u_div/PartRem[7][0] , \u_div/PartRem[6][0] , \u_div/PartRem[5][0] , 
        \u_div/PartRem[4][0] , \u_div/PartRem[3][0] , SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1}) );
  GSIM_DW_inc_2 \u_div/u_inc_QInc  ( .carry_in(n5), .a({n3, n3, n3, n4, 
        \u_div/QInv[59] , \u_div/QInv[58] , \u_div/QInv[57] , \u_div/QInv[56] , 
        \u_div/QInv[55] , \u_div/QInv[54] , \u_div/QInv[53] , \u_div/QInv[52] , 
        \u_div/QInv[51] , \u_div/QInv[50] , \u_div/QInv[49] , \u_div/QInv[48] , 
        \u_div/QInv[47] , \u_div/QInv[46] , \u_div/QInv[45] , \u_div/QInv[44] , 
        \u_div/QInv[43] , \u_div/QInv[42] , \u_div/QInv[41] , \u_div/QInv[40] , 
        \u_div/QInv[39] , \u_div/QInv[38] , \u_div/QInv[37] , \u_div/QInv[36] , 
        \u_div/QInv[35] , \u_div/QInv[34] , \u_div/QInv[33] , \u_div/QInv[32] , 
        \u_div/QInv[31] , \u_div/QInv[30] , \u_div/QInv[29] , \u_div/QInv[28] , 
        \u_div/QInv[27] , \u_div/QInv[26] , \u_div/QInv[25] , \u_div/QInv[24] , 
        \u_div/QInv[23] , \u_div/QInv[22] , \u_div/QInv[21] , \u_div/QInv[20] , 
        \u_div/QInv[19] , \u_div/QInv[18] , \u_div/QInv[17] , \u_div/QInv[16] , 
        \u_div/QInv[15] , \u_div/QInv[14] , \u_div/QInv[13] , \u_div/QInv[12] , 
        \u_div/QInv[11] , \u_div/QInv[10] , \u_div/QInv[9] , \u_div/QInv[8] , 
        \u_div/QInv[7] , \u_div/QInv[6] , \u_div/QInv[5] , \u_div/QInv[4] , 
        \u_div/QInv[3] , \u_div/QInv[2] , \u_div/QInv[1] , \u_div/QInv[0] }), 
        .sum(quotient) );
  ADDHXL \u_div/u_add_PartRem_2_4/U3  ( .A(\u_div/PartRem[5][4] ), .B(
        \u_div/u_add_PartRem_2_4/n3 ), .CO(\u_div/u_add_PartRem_2_4/n2 ), .S(
        \u_div/SumTmp[4][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_0  ( .A(\u_div/PartRem[3][0] ), .B(
        \u_div/PartRem[3][0] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/SumTmp[1][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_0  ( .A(\u_div/PartRem[21][0] ), .B(
        \u_div/PartRem[21][0] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/SumTmp[19][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_19_1  ( .A(\u_div/SumTmp[19][1] ), .B(
        \u_div/SumTmp[19][1] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_0  ( .A(\u_div/PartRem[26][0] ), .B(
        \u_div/PartRem[26][0] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/SumTmp[24][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_24_1  ( .A(\u_div/SumTmp[24][1] ), .B(
        \u_div/SumTmp[24][1] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_0  ( .A(\u_div/PartRem[31][0] ), .B(
        \u_div/PartRem[31][0] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/SumTmp[29][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_29_1  ( .A(\u_div/SumTmp[29][1] ), .B(
        \u_div/SumTmp[29][1] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_0  ( .A(\u_div/PartRem[36][0] ), .B(
        \u_div/PartRem[36][0] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/SumTmp[34][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_34_1  ( .A(\u_div/SumTmp[34][1] ), .B(
        \u_div/SumTmp[34][1] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_0  ( .A(\u_div/PartRem[41][0] ), .B(
        \u_div/PartRem[41][0] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/SumTmp[39][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_39_1  ( .A(\u_div/SumTmp[39][1] ), .B(
        \u_div/SumTmp[39][1] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_0  ( .A(\u_div/PartRem[46][0] ), .B(
        \u_div/PartRem[46][0] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/SumTmp[44][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_44_1  ( .A(\u_div/SumTmp[44][1] ), .B(
        \u_div/SumTmp[44][1] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_0  ( .A(\u_div/PartRem[51][0] ), .B(
        \u_div/PartRem[51][0] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/SumTmp[49][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_49_1  ( .A(\u_div/SumTmp[49][1] ), .B(
        \u_div/SumTmp[49][1] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_0  ( .A(\u_div/PartRem[56][0] ), .B(
        \u_div/PartRem[56][0] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/SumTmp[54][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_54_1  ( .A(\u_div/SumTmp[54][1] ), .B(
        \u_div/SumTmp[54][1] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_0  ( .A(\u_div/PartRem[5][0] ), .B(
        \u_div/PartRem[5][0] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/SumTmp[3][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_0  ( .A(\u_div/PartRem[6][0] ), .B(
        \u_div/PartRem[6][0] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/SumTmp[4][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_0  ( .A(\u_div/PartRem[8][0] ), .B(
        \u_div/PartRem[8][0] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/SumTmp[6][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_8_0  ( .A(\u_div/PartRem[9][0] ), .B(
        \u_div/PartRem[9][0] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/SumTmp[7][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_9_0  ( .A(\u_div/PartRem[10][0] ), .B(
        \u_div/PartRem[10][0] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/SumTmp[8][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_0  ( .A(\u_div/PartRem[11][0] ), .B(
        \u_div/PartRem[11][0] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/SumTmp[9][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_0  ( .A(\u_div/PartRem[13][0] ), .B(
        \u_div/PartRem[13][0] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/SumTmp[11][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_0  ( .A(\u_div/PartRem[14][0] ), .B(
        \u_div/PartRem[14][0] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/SumTmp[12][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_0  ( .A(\u_div/PartRem[16][0] ), .B(
        \u_div/PartRem[16][0] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/SumTmp[14][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_0  ( .A(\u_div/PartRem[15][0] ), .B(
        \u_div/PartRem[15][0] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/SumTmp[13][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_0  ( .A(\u_div/PartRem[17][0] ), .B(
        \u_div/PartRem[17][0] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/SumTmp[15][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_0  ( .A(\u_div/PartRem[18][0] ), .B(
        \u_div/PartRem[18][0] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/SumTmp[16][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_0  ( .A(\u_div/PartRem[19][0] ), .B(
        \u_div/PartRem[19][0] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/SumTmp[17][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_0  ( .A(\u_div/PartRem[22][0] ), .B(
        \u_div/PartRem[22][0] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/SumTmp[20][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_0  ( .A(\u_div/PartRem[23][0] ), .B(
        \u_div/PartRem[23][0] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/SumTmp[21][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_0  ( .A(\u_div/PartRem[24][0] ), .B(
        \u_div/PartRem[24][0] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/SumTmp[22][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_0  ( .A(\u_div/PartRem[27][0] ), .B(
        \u_div/PartRem[27][0] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/SumTmp[25][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_0  ( .A(\u_div/PartRem[28][0] ), .B(
        \u_div/PartRem[28][0] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/SumTmp[26][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_0  ( .A(\u_div/PartRem[29][0] ), .B(
        \u_div/PartRem[29][0] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/SumTmp[27][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_0  ( .A(\u_div/PartRem[32][0] ), .B(
        \u_div/PartRem[32][0] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/SumTmp[30][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_0  ( .A(\u_div/PartRem[34][0] ), .B(
        \u_div/PartRem[34][0] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/SumTmp[32][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_0  ( .A(\u_div/PartRem[37][0] ), .B(
        \u_div/PartRem[37][0] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/SumTmp[35][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_0  ( .A(\u_div/PartRem[38][0] ), .B(
        \u_div/PartRem[38][0] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/SumTmp[36][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_0  ( .A(\u_div/PartRem[39][0] ), .B(
        \u_div/PartRem[39][0] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/SumTmp[37][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_0  ( .A(\u_div/PartRem[42][0] ), .B(
        \u_div/PartRem[42][0] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/SumTmp[40][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_0  ( .A(\u_div/PartRem[43][0] ), .B(
        \u_div/PartRem[43][0] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/SumTmp[41][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_0  ( .A(\u_div/PartRem[44][0] ), .B(
        \u_div/PartRem[44][0] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/SumTmp[42][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_0  ( .A(\u_div/PartRem[47][0] ), .B(
        \u_div/PartRem[47][0] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/SumTmp[45][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_0  ( .A(\u_div/PartRem[48][0] ), .B(
        \u_div/PartRem[48][0] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/SumTmp[46][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_0  ( .A(\u_div/PartRem[49][0] ), .B(
        \u_div/PartRem[49][0] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/SumTmp[47][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_0  ( .A(\u_div/PartRem[52][0] ), .B(
        \u_div/PartRem[52][0] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/SumTmp[50][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_0  ( .A(\u_div/PartRem[53][0] ), .B(
        \u_div/PartRem[53][0] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/SumTmp[51][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_0  ( .A(\u_div/PartRem[54][0] ), .B(
        \u_div/PartRem[54][0] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/SumTmp[52][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_0  ( .A(\u_div/PartRem[57][0] ), .B(
        \u_div/PartRem[57][0] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/SumTmp[55][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_0  ( .A(\u_div/PartRem[58][0] ), .B(
        \u_div/PartRem[58][0] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/SumTmp[56][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_0  ( .A(\u_div/PartRem[59][0] ), .B(
        \u_div/PartRem[59][0] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/SumTmp[57][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_0  ( .A(\u_div/PartRem[4][0] ), .B(
        \u_div/PartRem[4][0] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/SumTmp[2][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_0  ( .A(\u_div/PartRem[7][0] ), .B(
        \u_div/PartRem[7][0] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/SumTmp[5][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_0  ( .A(\u_div/PartRem[12][0] ), .B(
        \u_div/PartRem[12][0] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/SumTmp[10][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_59_1  ( .A(\u_div/PartRem[61][0] ), .B(
        \u_div/PartRem[61][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_3  ( .A(\u_div/PartRem[4][3] ), .B(
        \u_div/SumTmp[3][3] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_3  ( .A(\u_div/PartRem[5][3] ), .B(
        \u_div/SumTmp[4][3] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_3  ( .A(\u_div/PartRem[8][3] ), .B(
        \u_div/SumTmp[7][3] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_8_3  ( .A(\u_div/PartRem[9][3] ), .B(
        \u_div/SumTmp[8][3] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_9_3  ( .A(\u_div/PartRem[10][3] ), .B(
        \u_div/SumTmp[9][3] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_3  ( .A(\u_div/PartRem[13][3] ), .B(
        \u_div/SumTmp[12][3] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_3  ( .A(\u_div/PartRem[7][3] ), .B(
        \u_div/SumTmp[6][3] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_3  ( .A(\u_div/PartRem[12][3] ), .B(
        \u_div/SumTmp[11][3] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_3  ( .A(\u_div/PartRem[15][3] ), .B(
        \u_div/SumTmp[14][3] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_1_3  ( .A(\u_div/PartRem[2][3] ), .B(
        \u_div/SumTmp[1][3] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_3  ( .A(\u_div/PartRem[3][3] ), .B(
        \u_div/SumTmp[2][3] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_3  ( .A(\u_div/PartRem[6][3] ), .B(
        \u_div/SumTmp[5][3] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_3  ( .A(\u_div/PartRem[17][3] ), .B(
        \u_div/SumTmp[16][3] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_3  ( .A(\u_div/PartRem[19][3] ), .B(
        \u_div/SumTmp[18][3] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_3  ( .A(\u_div/PartRem[21][3] ), .B(
        \u_div/SumTmp[20][3] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_3  ( .A(\u_div/PartRem[22][3] ), .B(
        \u_div/SumTmp[21][3] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_3  ( .A(\u_div/PartRem[24][3] ), .B(
        \u_div/SumTmp[23][3] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_3  ( .A(\u_div/PartRem[26][3] ), .B(
        \u_div/SumTmp[25][3] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_3  ( .A(\u_div/PartRem[27][3] ), .B(
        \u_div/SumTmp[26][3] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_3  ( .A(\u_div/PartRem[29][3] ), .B(
        \u_div/SumTmp[28][3] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_3  ( .A(\u_div/PartRem[31][3] ), .B(
        \u_div/SumTmp[30][3] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_3  ( .A(\u_div/PartRem[32][3] ), .B(
        \u_div/SumTmp[31][3] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_3  ( .A(\u_div/PartRem[34][3] ), .B(
        \u_div/SumTmp[33][3] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_3  ( .A(\u_div/PartRem[36][3] ), .B(
        \u_div/SumTmp[35][3] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_3  ( .A(\u_div/PartRem[37][3] ), .B(
        \u_div/SumTmp[36][3] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_3  ( .A(\u_div/PartRem[39][3] ), .B(
        \u_div/SumTmp[38][3] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_3  ( .A(\u_div/PartRem[41][3] ), .B(
        \u_div/SumTmp[40][3] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_3  ( .A(\u_div/PartRem[42][3] ), .B(
        \u_div/SumTmp[41][3] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_3  ( .A(\u_div/PartRem[44][3] ), .B(
        \u_div/SumTmp[43][3] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_3  ( .A(\u_div/PartRem[46][3] ), .B(
        \u_div/SumTmp[45][3] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_3  ( .A(\u_div/PartRem[47][3] ), .B(
        \u_div/SumTmp[46][3] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_3  ( .A(\u_div/PartRem[49][3] ), .B(
        \u_div/SumTmp[48][3] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_3  ( .A(\u_div/PartRem[51][3] ), .B(
        \u_div/SumTmp[50][3] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_3  ( .A(\u_div/PartRem[52][3] ), .B(
        \u_div/SumTmp[51][3] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_3  ( .A(\u_div/PartRem[54][3] ), .B(
        \u_div/SumTmp[53][3] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_3  ( .A(\u_div/PartRem[56][3] ), .B(
        \u_div/SumTmp[55][3] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_3  ( .A(\u_div/PartRem[57][3] ), .B(
        \u_div/SumTmp[56][3] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_3  ( .A(\u_div/PartRem[59][3] ), .B(
        \u_div/SumTmp[58][3] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_3  ( .A(\u_div/PartRem[11][3] ), .B(
        \u_div/SumTmp[10][3] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_3  ( .A(\u_div/PartRem[14][3] ), .B(
        \u_div/SumTmp[13][3] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_3  ( .A(\u_div/PartRem[23][3] ), .B(
        \u_div/SumTmp[22][3] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_3  ( .A(\u_div/PartRem[28][3] ), .B(
        \u_div/SumTmp[27][3] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_3  ( .A(\u_div/PartRem[38][3] ), .B(
        \u_div/SumTmp[37][3] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_3  ( .A(\u_div/PartRem[43][3] ), .B(
        \u_div/SumTmp[42][3] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_3  ( .A(\u_div/PartRem[48][3] ), .B(
        \u_div/SumTmp[47][3] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_3  ( .A(\u_div/PartRem[53][3] ), .B(
        \u_div/SumTmp[52][3] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_3  ( .A(\u_div/PartRem[58][3] ), .B(
        \u_div/SumTmp[57][3] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_3  ( .A(\u_div/PartRem[16][3] ), .B(
        \u_div/SumTmp[15][3] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_3  ( .A(\u_div/PartRem[18][3] ), .B(
        \u_div/SumTmp[17][3] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_3  ( .A(\u_div/PartRem[33][3] ), .B(
        \u_div/SumTmp[32][3] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/SumTmp[1][2] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_3_1  ( .A(\u_div/SumTmp[3][1] ), .B(
        \u_div/SumTmp[3][1] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_4_1  ( .A(\u_div/SumTmp[4][1] ), .B(
        \u_div/SumTmp[4][1] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_6_1  ( .A(\u_div/SumTmp[6][1] ), .B(
        \u_div/SumTmp[6][1] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_7_1  ( .A(\u_div/SumTmp[7][1] ), .B(
        \u_div/SumTmp[7][1] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_8_1  ( .A(\u_div/SumTmp[8][1] ), .B(
        \u_div/SumTmp[8][1] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_9_1  ( .A(\u_div/SumTmp[9][1] ), .B(
        \u_div/SumTmp[9][1] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_11_1  ( .A(\u_div/SumTmp[11][1] ), .B(
        \u_div/SumTmp[11][1] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_14_1  ( .A(\u_div/SumTmp[14][1] ), .B(
        \u_div/SumTmp[14][1] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_12_1  ( .A(\u_div/SumTmp[12][1] ), .B(
        \u_div/SumTmp[12][1] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_5_1  ( .A(\u_div/SumTmp[5][1] ), .B(
        \u_div/SumTmp[5][1] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_10_1  ( .A(\u_div/SumTmp[10][1] ), .B(
        \u_div/SumTmp[10][1] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_17_1  ( .A(\u_div/SumTmp[17][1] ), .B(
        \u_div/SumTmp[17][1] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_16_1  ( .A(\u_div/SumTmp[16][1] ), .B(
        \u_div/SumTmp[16][1] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_15_1  ( .A(\u_div/SumTmp[15][1] ), .B(
        \u_div/SumTmp[15][1] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_13_1  ( .A(\u_div/SumTmp[13][1] ), .B(
        \u_div/SumTmp[13][1] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_18_1  ( .A(\u_div/SumTmp[18][1] ), .B(
        \u_div/SumTmp[18][1] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_0  ( .A(\u_div/PartRem[20][0] ), .B(
        \u_div/PartRem[20][0] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/SumTmp[18][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_22_1  ( .A(\u_div/SumTmp[22][1] ), .B(
        \u_div/SumTmp[22][1] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_21_1  ( .A(\u_div/SumTmp[21][1] ), .B(
        \u_div/SumTmp[21][1] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_20_1  ( .A(\u_div/SumTmp[20][1] ), .B(
        \u_div/SumTmp[20][1] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_23_1  ( .A(\u_div/SumTmp[23][1] ), .B(
        \u_div/SumTmp[23][1] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_0  ( .A(\u_div/PartRem[25][0] ), .B(
        \u_div/PartRem[25][0] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/SumTmp[23][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_25_1  ( .A(\u_div/SumTmp[25][1] ), .B(
        \u_div/SumTmp[25][1] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_26_1  ( .A(\u_div/SumTmp[26][1] ), .B(
        \u_div/SumTmp[26][1] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_27_1  ( .A(\u_div/SumTmp[27][1] ), .B(
        \u_div/SumTmp[27][1] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_28_1  ( .A(\u_div/SumTmp[28][1] ), .B(
        \u_div/SumTmp[28][1] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_0  ( .A(\u_div/PartRem[30][0] ), .B(
        \u_div/PartRem[30][0] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/SumTmp[28][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_30_1  ( .A(\u_div/SumTmp[30][1] ), .B(
        \u_div/SumTmp[30][1] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_31_1  ( .A(\u_div/SumTmp[31][1] ), .B(
        \u_div/SumTmp[31][1] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_33_1  ( .A(\u_div/SumTmp[33][1] ), .B(
        \u_div/SumTmp[33][1] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_0  ( .A(\u_div/PartRem[35][0] ), .B(
        \u_div/PartRem[35][0] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/SumTmp[33][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_35_1  ( .A(\u_div/SumTmp[35][1] ), .B(
        \u_div/SumTmp[35][1] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_36_1  ( .A(\u_div/SumTmp[36][1] ), .B(
        \u_div/SumTmp[36][1] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_37_1  ( .A(\u_div/SumTmp[37][1] ), .B(
        \u_div/SumTmp[37][1] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_38_1  ( .A(\u_div/SumTmp[38][1] ), .B(
        \u_div/SumTmp[38][1] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_0  ( .A(\u_div/PartRem[40][0] ), .B(
        \u_div/PartRem[40][0] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/SumTmp[38][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_40_1  ( .A(\u_div/SumTmp[40][1] ), .B(
        \u_div/SumTmp[40][1] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_41_1  ( .A(\u_div/SumTmp[41][1] ), .B(
        \u_div/SumTmp[41][1] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_42_1  ( .A(\u_div/SumTmp[42][1] ), .B(
        \u_div/SumTmp[42][1] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_43_1  ( .A(\u_div/SumTmp[43][1] ), .B(
        \u_div/SumTmp[43][1] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_0  ( .A(\u_div/PartRem[45][0] ), .B(
        \u_div/PartRem[45][0] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/SumTmp[43][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_45_1  ( .A(\u_div/SumTmp[45][1] ), .B(
        \u_div/SumTmp[45][1] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_46_1  ( .A(\u_div/SumTmp[46][1] ), .B(
        \u_div/SumTmp[46][1] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_47_1  ( .A(\u_div/SumTmp[47][1] ), .B(
        \u_div/SumTmp[47][1] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_48_1  ( .A(\u_div/SumTmp[48][1] ), .B(
        \u_div/SumTmp[48][1] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_0  ( .A(\u_div/PartRem[50][0] ), .B(
        \u_div/PartRem[50][0] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/SumTmp[48][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_51_1  ( .A(\u_div/SumTmp[51][1] ), .B(
        \u_div/SumTmp[51][1] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_50_1  ( .A(\u_div/SumTmp[50][1] ), .B(
        \u_div/SumTmp[50][1] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_52_1  ( .A(\u_div/SumTmp[52][1] ), .B(
        \u_div/SumTmp[52][1] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_53_1  ( .A(\u_div/SumTmp[53][1] ), .B(
        \u_div/SumTmp[53][1] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_0  ( .A(\u_div/PartRem[55][0] ), .B(
        \u_div/PartRem[55][0] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/SumTmp[53][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_55_1  ( .A(\u_div/SumTmp[55][1] ), .B(
        \u_div/SumTmp[55][1] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_56_1  ( .A(\u_div/SumTmp[56][1] ), .B(
        \u_div/SumTmp[56][1] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_57_1  ( .A(\u_div/SumTmp[57][1] ), .B(
        \u_div/SumTmp[57][1] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_58_1  ( .A(\u_div/SumTmp[58][1] ), .B(
        \u_div/SumTmp[58][1] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_0  ( .A(\u_div/PartRem[60][0] ), .B(
        \u_div/PartRem[60][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/SumTmp[58][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_2_1  ( .A(\u_div/SumTmp[2][1] ), .B(
        \u_div/SumTmp[2][1] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_3  ( .A(\u_div/PartRem[20][3] ), .B(
        \u_div/SumTmp[19][3] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_3  ( .A(\u_div/PartRem[25][3] ), .B(
        \u_div/SumTmp[24][3] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_3  ( .A(\u_div/PartRem[30][3] ), .B(
        \u_div/SumTmp[29][3] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_3  ( .A(\u_div/PartRem[35][3] ), .B(
        \u_div/SumTmp[34][3] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_3  ( .A(\u_div/PartRem[40][3] ), .B(
        \u_div/SumTmp[39][3] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_3  ( .A(\u_div/PartRem[45][3] ), .B(
        \u_div/SumTmp[44][3] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_3  ( .A(\u_div/PartRem[50][3] ), .B(
        \u_div/SumTmp[49][3] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_3  ( .A(\u_div/PartRem[55][3] ), .B(
        \u_div/SumTmp[54][3] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_3  ( .A(\u_div/PartRem[63][0] ), .B(
        \u_div/SumTmp[59][3] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_1_4  ( .A(\u_div/PartRem[2][4] ), .B(
        \u_div/SumTmp[1][4] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_4  ( .A(\u_div/PartRem[21][4] ), .B(
        \u_div/SumTmp[20][4] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_4  ( .A(\u_div/PartRem[26][4] ), .B(
        \u_div/SumTmp[25][4] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_4  ( .A(\u_div/PartRem[31][4] ), .B(
        \u_div/SumTmp[30][4] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_4  ( .A(\u_div/PartRem[36][4] ), .B(
        \u_div/SumTmp[35][4] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_4  ( .A(\u_div/PartRem[41][4] ), .B(
        \u_div/SumTmp[40][4] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_4  ( .A(\u_div/PartRem[46][4] ), .B(
        \u_div/SumTmp[45][4] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_4  ( .A(\u_div/PartRem[51][4] ), .B(
        \u_div/SumTmp[50][4] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_4  ( .A(\u_div/PartRem[56][4] ), .B(
        \u_div/SumTmp[55][4] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_4  ( .A(\u_div/PartRem[3][4] ), .B(
        \u_div/SumTmp[2][4] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_4  ( .A(\u_div/PartRem[4][4] ), .B(
        \u_div/SumTmp[3][4] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_4  ( .A(\u_div/PartRem[5][4] ), .B(
        \u_div/SumTmp[4][4] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_4  ( .A(\u_div/PartRem[6][4] ), .B(
        \u_div/SumTmp[5][4] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_4  ( .A(\u_div/PartRem[8][4] ), .B(
        \u_div/SumTmp[7][4] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_8_4  ( .A(\u_div/PartRem[9][4] ), .B(
        \u_div/SumTmp[8][4] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_9_4  ( .A(\u_div/PartRem[10][4] ), .B(
        \u_div/SumTmp[9][4] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_4  ( .A(\u_div/PartRem[11][4] ), .B(
        \u_div/SumTmp[10][4] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_4  ( .A(\u_div/PartRem[13][4] ), .B(
        \u_div/SumTmp[12][4] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_4  ( .A(\u_div/PartRem[14][4] ), .B(
        \u_div/SumTmp[13][4] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_4  ( .A(\u_div/PartRem[16][4] ), .B(
        \u_div/SumTmp[15][4] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_4  ( .A(\u_div/PartRem[7][4] ), .B(
        \u_div/SumTmp[6][4] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_4  ( .A(\u_div/PartRem[12][4] ), .B(
        \u_div/SumTmp[11][4] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_4  ( .A(\u_div/PartRem[15][4] ), .B(
        \u_div/SumTmp[14][4] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_4  ( .A(\u_div/PartRem[18][4] ), .B(
        \u_div/SumTmp[17][4] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_4  ( .A(\u_div/PartRem[19][4] ), .B(
        \u_div/SumTmp[18][4] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_4  ( .A(\u_div/PartRem[17][4] ), .B(
        \u_div/SumTmp[16][4] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_4  ( .A(\u_div/PartRem[20][4] ), .B(
        \u_div/SumTmp[19][4] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_4  ( .A(\u_div/PartRem[23][4] ), .B(
        \u_div/SumTmp[22][4] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_4  ( .A(\u_div/PartRem[22][4] ), .B(
        \u_div/SumTmp[21][4] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_4  ( .A(\u_div/PartRem[24][4] ), .B(
        \u_div/SumTmp[23][4] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_4  ( .A(\u_div/PartRem[25][4] ), .B(
        \u_div/SumTmp[24][4] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_4  ( .A(\u_div/PartRem[29][4] ), .B(
        \u_div/SumTmp[28][4] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_4  ( .A(\u_div/PartRem[27][4] ), .B(
        \u_div/SumTmp[26][4] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_4  ( .A(\u_div/PartRem[28][4] ), .B(
        \u_div/SumTmp[27][4] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_4  ( .A(\u_div/PartRem[30][4] ), .B(
        \u_div/SumTmp[29][4] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_4  ( .A(\u_div/PartRem[34][4] ), .B(
        \u_div/SumTmp[33][4] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_4  ( .A(\u_div/PartRem[32][4] ), .B(
        \u_div/SumTmp[31][4] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_4  ( .A(\u_div/PartRem[35][4] ), .B(
        \u_div/SumTmp[34][4] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_4  ( .A(\u_div/PartRem[37][4] ), .B(
        \u_div/SumTmp[36][4] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_4  ( .A(\u_div/PartRem[39][4] ), .B(
        \u_div/SumTmp[38][4] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_4  ( .A(\u_div/PartRem[38][4] ), .B(
        \u_div/SumTmp[37][4] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_4  ( .A(\u_div/PartRem[40][4] ), .B(
        \u_div/SumTmp[39][4] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_4  ( .A(\u_div/PartRem[44][4] ), .B(
        \u_div/SumTmp[43][4] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_4  ( .A(\u_div/PartRem[42][4] ), .B(
        \u_div/SumTmp[41][4] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_4  ( .A(\u_div/PartRem[43][4] ), .B(
        \u_div/SumTmp[42][4] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_4  ( .A(\u_div/PartRem[47][4] ), .B(
        \u_div/SumTmp[46][4] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_4  ( .A(\u_div/PartRem[50][4] ), .B(
        \u_div/SumTmp[49][4] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_4  ( .A(\u_div/PartRem[45][4] ), .B(
        \u_div/SumTmp[44][4] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_4  ( .A(\u_div/PartRem[52][4] ), .B(
        \u_div/SumTmp[51][4] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_4  ( .A(\u_div/PartRem[49][4] ), .B(
        \u_div/SumTmp[48][4] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_4  ( .A(\u_div/PartRem[48][4] ), .B(
        \u_div/SumTmp[47][4] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_4  ( .A(\u_div/PartRem[55][4] ), .B(
        \u_div/SumTmp[54][4] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_4  ( .A(\u_div/PartRem[53][4] ), .B(
        \u_div/SumTmp[52][4] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_4  ( .A(\u_div/PartRem[54][4] ), .B(
        \u_div/SumTmp[53][4] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_4  ( .A(\u_div/PartRem[58][4] ), .B(
        \u_div/SumTmp[57][4] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_4  ( .A(\u_div/PartRem[57][4] ), .B(
        \u_div/SumTmp[56][4] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_4  ( .A(\u_div/PartRem[59][4] ), .B(
        \u_div/SumTmp[58][4] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_4  ( .A(\u_div/PartRem[64][0] ), .B(
        \u_div/SumTmp[59][4] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_32_4  ( .A(\u_div/PartRem[33][4] ), .B(
        \u_div/SumTmp[32][4] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_32_1  ( .A(\u_div/SumTmp[32][1] ), .B(
        \u_div/SumTmp[32][1] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_32_0  ( .A(\u_div/PartRem[33][0] ), .B(
        \u_div/PartRem[33][0] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/SumTmp[31][1] ) );
  OR2X8 U1 ( .A(\u_div/PartRem[48][5] ), .B(\u_div/u_add_PartRem_2_47/n2 ), 
        .Y(\u_div/CryTmp[47][6] ) );
  ADDHX2 U2 ( .A(\u_div/PartRem[48][4] ), .B(\u_div/u_add_PartRem_2_47/n3 ), 
        .CO(\u_div/u_add_PartRem_2_47/n2 ), .S(\u_div/SumTmp[47][4] ) );
  MXI2X2 U3 ( .A(\u_div/SumTmp[32][2] ), .B(\u_div/PartRem[33][2] ), .S0(
        \u_div/CryTmp[32][6] ), .Y(\u_div/PartRem[32][3] ) );
  OR2X6 U4 ( .A(\u_div/PartRem[14][5] ), .B(\u_div/u_add_PartRem_2_13/n2 ), 
        .Y(\u_div/CryTmp[13][6] ) );
  OR2X6 U5 ( .A(\u_div/PartRem[16][5] ), .B(\u_div/u_add_PartRem_2_15/n2 ), 
        .Y(\u_div/CryTmp[15][6] ) );
  OR2X6 U6 ( .A(\u_div/PartRem[18][5] ), .B(\u_div/u_add_PartRem_2_17/n2 ), 
        .Y(\u_div/CryTmp[17][6] ) );
  OR2X6 U7 ( .A(\u_div/PartRem[23][5] ), .B(\u_div/u_add_PartRem_2_22/n2 ), 
        .Y(\u_div/CryTmp[22][6] ) );
  OR2X6 U8 ( .A(\u_div/PartRem[28][5] ), .B(\u_div/u_add_PartRem_2_27/n2 ), 
        .Y(\u_div/CryTmp[27][6] ) );
  OR2X6 U9 ( .A(\u_div/PartRem[38][5] ), .B(\u_div/u_add_PartRem_2_37/n2 ), 
        .Y(\u_div/CryTmp[37][6] ) );
  OR2X6 U10 ( .A(\u_div/PartRem[43][5] ), .B(\u_div/u_add_PartRem_2_42/n2 ), 
        .Y(\u_div/CryTmp[42][6] ) );
  OR2X6 U11 ( .A(\u_div/PartRem[59][5] ), .B(\u_div/u_add_PartRem_2_58/n2 ), 
        .Y(\u_div/CryTmp[58][6] ) );
  ADDHX2 U12 ( .A(\u_div/PartRem[43][4] ), .B(\u_div/u_add_PartRem_2_42/n3 ), 
        .CO(\u_div/u_add_PartRem_2_42/n2 ), .S(\u_div/SumTmp[42][4] ) );
  ADDHX2 U13 ( .A(\u_div/PartRem[38][4] ), .B(\u_div/u_add_PartRem_2_37/n3 ), 
        .CO(\u_div/u_add_PartRem_2_37/n2 ), .S(\u_div/SumTmp[37][4] ) );
  ADDHX2 U14 ( .A(\u_div/PartRem[28][4] ), .B(\u_div/u_add_PartRem_2_27/n3 ), 
        .CO(\u_div/u_add_PartRem_2_27/n2 ), .S(\u_div/SumTmp[27][4] ) );
  ADDHX2 U15 ( .A(\u_div/PartRem[23][4] ), .B(\u_div/u_add_PartRem_2_22/n3 ), 
        .CO(\u_div/u_add_PartRem_2_22/n2 ), .S(\u_div/SumTmp[22][4] ) );
  ADDHX2 U16 ( .A(\u_div/PartRem[16][4] ), .B(\u_div/u_add_PartRem_2_15/n3 ), 
        .CO(\u_div/u_add_PartRem_2_15/n2 ), .S(\u_div/SumTmp[15][4] ) );
  OR2X8 U17 ( .A(\u_div/PartRem[58][5] ), .B(\u_div/u_add_PartRem_2_57/n2 ), 
        .Y(\u_div/CryTmp[57][6] ) );
  ADDHX2 U18 ( .A(\u_div/PartRem[58][4] ), .B(\u_div/u_add_PartRem_2_57/n3 ), 
        .CO(\u_div/u_add_PartRem_2_57/n2 ), .S(\u_div/SumTmp[57][4] ) );
  XOR2XL U19 ( .A(\u_div/CryTmp[32][6] ), .B(n3), .Y(\u_div/QInv[32] ) );
  OR2X6 U20 ( .A(\u_div/PartRem[33][5] ), .B(\u_div/u_add_PartRem_2_32/n2 ), 
        .Y(\u_div/CryTmp[32][6] ) );
  ADDHX2 U21 ( .A(\u_div/PartRem[18][4] ), .B(\u_div/u_add_PartRem_2_17/n3 ), 
        .CO(\u_div/u_add_PartRem_2_17/n2 ), .S(\u_div/SumTmp[17][4] ) );
  ADDHX2 U22 ( .A(\u_div/PartRem[14][4] ), .B(\u_div/u_add_PartRem_2_13/n3 ), 
        .CO(\u_div/u_add_PartRem_2_13/n2 ), .S(\u_div/SumTmp[13][4] ) );
  ADDHX2 U23 ( .A(\u_div/PartRem[59][4] ), .B(\u_div/u_add_PartRem_2_58/n3 ), 
        .CO(\u_div/u_add_PartRem_2_58/n2 ), .S(\u_div/SumTmp[58][4] ) );
  NOR2X4 U24 ( .A(\u_div/PartRem[63][0] ), .B(\u_div/PartRem[62][0] ), .Y(n8)
         );
  OR2X1 U25 ( .A(\u_div/PartRem[55][5] ), .B(\u_div/u_add_PartRem_2_54/n2 ), 
        .Y(\u_div/CryTmp[54][6] ) );
  OR2X1 U26 ( .A(\u_div/PartRem[45][5] ), .B(\u_div/u_add_PartRem_2_44/n2 ), 
        .Y(\u_div/CryTmp[44][6] ) );
  OR2X1 U27 ( .A(\u_div/PartRem[50][5] ), .B(\u_div/u_add_PartRem_2_49/n2 ), 
        .Y(\u_div/CryTmp[49][6] ) );
  OR2X1 U28 ( .A(\u_div/PartRem[40][5] ), .B(\u_div/u_add_PartRem_2_39/n2 ), 
        .Y(\u_div/CryTmp[39][6] ) );
  OR2X1 U29 ( .A(\u_div/PartRem[35][5] ), .B(\u_div/u_add_PartRem_2_34/n2 ), 
        .Y(\u_div/CryTmp[34][6] ) );
  OR2X1 U30 ( .A(\u_div/PartRem[30][5] ), .B(\u_div/u_add_PartRem_2_29/n2 ), 
        .Y(\u_div/CryTmp[29][6] ) );
  OR2X1 U31 ( .A(\u_div/PartRem[25][5] ), .B(\u_div/u_add_PartRem_2_24/n2 ), 
        .Y(\u_div/CryTmp[24][6] ) );
  OR2X1 U32 ( .A(\u_div/PartRem[20][5] ), .B(\u_div/u_add_PartRem_2_19/n2 ), 
        .Y(\u_div/CryTmp[19][6] ) );
  ADDHXL U33 ( .A(\u_div/PartRem[55][4] ), .B(\u_div/u_add_PartRem_2_54/n3 ), 
        .CO(\u_div/u_add_PartRem_2_54/n2 ), .S(\u_div/SumTmp[54][4] ) );
  ADDHXL U34 ( .A(\u_div/PartRem[31][4] ), .B(\u_div/u_add_PartRem_2_30/n3 ), 
        .CO(\u_div/u_add_PartRem_2_30/n2 ), .S(\u_div/SumTmp[30][4] ) );
  ADDHXL U35 ( .A(\u_div/PartRem[56][4] ), .B(\u_div/u_add_PartRem_2_55/n3 ), 
        .CO(\u_div/u_add_PartRem_2_55/n2 ), .S(\u_div/SumTmp[55][4] ) );
  ADDHXL U36 ( .A(\u_div/PartRem[53][4] ), .B(\u_div/u_add_PartRem_2_52/n3 ), 
        .CO(\u_div/u_add_PartRem_2_52/n2 ), .S(\u_div/SumTmp[52][4] ) );
  ADDHXL U37 ( .A(\u_div/PartRem[51][4] ), .B(\u_div/u_add_PartRem_2_50/n3 ), 
        .CO(\u_div/u_add_PartRem_2_50/n2 ), .S(\u_div/SumTmp[50][4] ) );
  ADDHXL U38 ( .A(\u_div/PartRem[50][4] ), .B(\u_div/u_add_PartRem_2_49/n3 ), 
        .CO(\u_div/u_add_PartRem_2_49/n2 ), .S(\u_div/SumTmp[49][4] ) );
  ADDHXL U39 ( .A(\u_div/PartRem[46][4] ), .B(\u_div/u_add_PartRem_2_45/n3 ), 
        .CO(\u_div/u_add_PartRem_2_45/n2 ), .S(\u_div/SumTmp[45][4] ) );
  ADDHXL U40 ( .A(\u_div/PartRem[45][4] ), .B(\u_div/u_add_PartRem_2_44/n3 ), 
        .CO(\u_div/u_add_PartRem_2_44/n2 ), .S(\u_div/SumTmp[44][4] ) );
  ADDHXL U41 ( .A(\u_div/PartRem[41][4] ), .B(\u_div/u_add_PartRem_2_40/n3 ), 
        .CO(\u_div/u_add_PartRem_2_40/n2 ), .S(\u_div/SumTmp[40][4] ) );
  ADDHXL U42 ( .A(\u_div/PartRem[40][4] ), .B(\u_div/u_add_PartRem_2_39/n3 ), 
        .CO(\u_div/u_add_PartRem_2_39/n2 ), .S(\u_div/SumTmp[39][4] ) );
  ADDHXL U43 ( .A(\u_div/PartRem[36][4] ), .B(\u_div/u_add_PartRem_2_35/n3 ), 
        .CO(\u_div/u_add_PartRem_2_35/n2 ), .S(\u_div/SumTmp[35][4] ) );
  ADDHXL U44 ( .A(\u_div/PartRem[35][4] ), .B(\u_div/u_add_PartRem_2_34/n3 ), 
        .CO(\u_div/u_add_PartRem_2_34/n2 ), .S(\u_div/SumTmp[34][4] ) );
  ADDHXL U45 ( .A(\u_div/PartRem[33][4] ), .B(\u_div/u_add_PartRem_2_32/n3 ), 
        .CO(\u_div/u_add_PartRem_2_32/n2 ), .S(\u_div/SumTmp[32][4] ) );
  ADDHXL U46 ( .A(\u_div/PartRem[30][4] ), .B(\u_div/u_add_PartRem_2_29/n3 ), 
        .CO(\u_div/u_add_PartRem_2_29/n2 ), .S(\u_div/SumTmp[29][4] ) );
  ADDHXL U47 ( .A(\u_div/PartRem[26][4] ), .B(\u_div/u_add_PartRem_2_25/n3 ), 
        .CO(\u_div/u_add_PartRem_2_25/n2 ), .S(\u_div/SumTmp[25][4] ) );
  ADDHXL U48 ( .A(\u_div/PartRem[25][4] ), .B(\u_div/u_add_PartRem_2_24/n3 ), 
        .CO(\u_div/u_add_PartRem_2_24/n2 ), .S(\u_div/SumTmp[24][4] ) );
  ADDHXL U49 ( .A(\u_div/PartRem[21][4] ), .B(\u_div/u_add_PartRem_2_20/n3 ), 
        .CO(\u_div/u_add_PartRem_2_20/n2 ), .S(\u_div/SumTmp[20][4] ) );
  ADDHXL U50 ( .A(\u_div/PartRem[20][4] ), .B(\u_div/u_add_PartRem_2_19/n3 ), 
        .CO(\u_div/u_add_PartRem_2_19/n2 ), .S(\u_div/SumTmp[19][4] ) );
  ADDHXL U51 ( .A(\u_div/PartRem[12][4] ), .B(\u_div/u_add_PartRem_2_11/n3 ), 
        .CO(\u_div/u_add_PartRem_2_11/n2 ), .S(\u_div/SumTmp[11][4] ) );
  ADDHXL U52 ( .A(\u_div/PartRem[11][4] ), .B(\u_div/u_add_PartRem_2_10/n3 ), 
        .CO(\u_div/u_add_PartRem_2_10/n2 ), .S(\u_div/SumTmp[10][4] ) );
  ADDHXL U53 ( .A(\u_div/PartRem[10][4] ), .B(\u_div/u_add_PartRem_2_9/n3 ), 
        .CO(\u_div/u_add_PartRem_2_9/n2 ), .S(\u_div/SumTmp[9][4] ) );
  ADDHXL U54 ( .A(\u_div/PartRem[9][4] ), .B(\u_div/u_add_PartRem_2_8/n3 ), 
        .CO(\u_div/u_add_PartRem_2_8/n2 ), .S(\u_div/SumTmp[8][4] ) );
  ADDHXL U55 ( .A(\u_div/PartRem[8][4] ), .B(\u_div/u_add_PartRem_2_7/n3 ), 
        .CO(\u_div/u_add_PartRem_2_7/n2 ), .S(\u_div/SumTmp[7][4] ) );
  ADDHXL U56 ( .A(\u_div/PartRem[7][4] ), .B(\u_div/u_add_PartRem_2_6/n3 ), 
        .CO(\u_div/u_add_PartRem_2_6/n2 ), .S(\u_div/SumTmp[6][4] ) );
  ADDHXL U57 ( .A(\u_div/PartRem[6][4] ), .B(\u_div/u_add_PartRem_2_5/n3 ), 
        .CO(\u_div/u_add_PartRem_2_5/n2 ), .S(\u_div/SumTmp[5][4] ) );
  ADDHXL U58 ( .A(\u_div/PartRem[4][4] ), .B(\u_div/u_add_PartRem_2_3/n3 ), 
        .CO(\u_div/u_add_PartRem_2_3/n2 ), .S(\u_div/SumTmp[3][4] ) );
  ADDHXL U59 ( .A(\u_div/PartRem[3][4] ), .B(\u_div/u_add_PartRem_2_2/n3 ), 
        .CO(\u_div/u_add_PartRem_2_2/n2 ), .S(\u_div/SumTmp[2][4] ) );
  ADDHXL U60 ( .A(\u_div/PartRem[2][4] ), .B(\u_div/u_add_PartRem_2_1/n3 ), 
        .CO(\u_div/u_add_PartRem_2_1/n2 ), .S(\u_div/SumTmp[1][4] ) );
  ADDHXL U61 ( .A(\u_div/PartRem[54][4] ), .B(\u_div/u_add_PartRem_2_53/n3 ), 
        .CO(\u_div/u_add_PartRem_2_53/n2 ), .S(\u_div/SumTmp[53][4] ) );
  ADDHXL U62 ( .A(\u_div/PartRem[49][4] ), .B(\u_div/u_add_PartRem_2_48/n3 ), 
        .CO(\u_div/u_add_PartRem_2_48/n2 ), .S(\u_div/SumTmp[48][4] ) );
  ADDHXL U63 ( .A(\u_div/PartRem[44][4] ), .B(\u_div/u_add_PartRem_2_43/n3 ), 
        .CO(\u_div/u_add_PartRem_2_43/n2 ), .S(\u_div/SumTmp[43][4] ) );
  ADDHXL U64 ( .A(\u_div/PartRem[39][4] ), .B(\u_div/u_add_PartRem_2_38/n3 ), 
        .CO(\u_div/u_add_PartRem_2_38/n2 ), .S(\u_div/SumTmp[38][4] ) );
  ADDHXL U65 ( .A(\u_div/PartRem[34][4] ), .B(\u_div/u_add_PartRem_2_33/n3 ), 
        .CO(\u_div/u_add_PartRem_2_33/n2 ), .S(\u_div/SumTmp[33][4] ) );
  ADDHXL U66 ( .A(\u_div/PartRem[29][4] ), .B(\u_div/u_add_PartRem_2_28/n3 ), 
        .CO(\u_div/u_add_PartRem_2_28/n2 ), .S(\u_div/SumTmp[28][4] ) );
  ADDHXL U67 ( .A(\u_div/PartRem[24][4] ), .B(\u_div/u_add_PartRem_2_23/n3 ), 
        .CO(\u_div/u_add_PartRem_2_23/n2 ), .S(\u_div/SumTmp[23][4] ) );
  ADDHXL U68 ( .A(\u_div/PartRem[19][4] ), .B(\u_div/u_add_PartRem_2_18/n3 ), 
        .CO(\u_div/u_add_PartRem_2_18/n2 ), .S(\u_div/SumTmp[18][4] ) );
  ADDHXL U69 ( .A(\u_div/PartRem[27][4] ), .B(\u_div/u_add_PartRem_2_26/n3 ), 
        .CO(\u_div/u_add_PartRem_2_26/n2 ), .S(\u_div/SumTmp[26][4] ) );
  ADDHXL U70 ( .A(\u_div/PartRem[32][4] ), .B(\u_div/u_add_PartRem_2_31/n3 ), 
        .CO(\u_div/u_add_PartRem_2_31/n2 ), .S(\u_div/SumTmp[31][4] ) );
  ADDHXL U71 ( .A(\u_div/PartRem[17][4] ), .B(\u_div/u_add_PartRem_2_16/n3 ), 
        .CO(\u_div/u_add_PartRem_2_16/n2 ), .S(\u_div/SumTmp[16][4] ) );
  ADDHXL U72 ( .A(\u_div/PartRem[37][4] ), .B(\u_div/u_add_PartRem_2_36/n3 ), 
        .CO(\u_div/u_add_PartRem_2_36/n2 ), .S(\u_div/SumTmp[36][4] ) );
  ADDHXL U73 ( .A(\u_div/PartRem[22][4] ), .B(\u_div/u_add_PartRem_2_21/n3 ), 
        .CO(\u_div/u_add_PartRem_2_21/n2 ), .S(\u_div/SumTmp[21][4] ) );
  ADDHXL U74 ( .A(\u_div/PartRem[42][4] ), .B(\u_div/u_add_PartRem_2_41/n3 ), 
        .CO(\u_div/u_add_PartRem_2_41/n2 ), .S(\u_div/SumTmp[41][4] ) );
  ADDHXL U75 ( .A(\u_div/PartRem[57][4] ), .B(\u_div/u_add_PartRem_2_56/n3 ), 
        .CO(\u_div/u_add_PartRem_2_56/n2 ), .S(\u_div/SumTmp[56][4] ) );
  ADDHXL U76 ( .A(\u_div/PartRem[15][4] ), .B(\u_div/u_add_PartRem_2_14/n3 ), 
        .CO(\u_div/u_add_PartRem_2_14/n2 ), .S(\u_div/SumTmp[14][4] ) );
  ADDHXL U77 ( .A(\u_div/PartRem[47][4] ), .B(\u_div/u_add_PartRem_2_46/n3 ), 
        .CO(\u_div/u_add_PartRem_2_46/n2 ), .S(\u_div/SumTmp[46][4] ) );
  ADDHXL U78 ( .A(\u_div/PartRem[13][4] ), .B(\u_div/u_add_PartRem_2_12/n3 ), 
        .CO(\u_div/u_add_PartRem_2_12/n2 ), .S(\u_div/SumTmp[12][4] ) );
  ADDHXL U79 ( .A(\u_div/PartRem[52][4] ), .B(\u_div/u_add_PartRem_2_51/n3 ), 
        .CO(\u_div/u_add_PartRem_2_51/n2 ), .S(\u_div/SumTmp[51][4] ) );
  NOR2BX4 U80 ( .AN(\u_div/PartRem[64][0] ), .B(n8), .Y(\u_div/CryTmp[59][6] )
         );
  AO21X4 U81 ( .A0(\u_div/PartRem[1][4] ), .A1(n6), .B0(\u_div/PartRem[1][5] ), 
        .Y(\u_div/CryTmp[0][6] ) );
  MXI2X2 U82 ( .A(\u_div/SumTmp[17][2] ), .B(\u_div/PartRem[18][2] ), .S0(
        \u_div/CryTmp[17][6] ), .Y(\u_div/PartRem[17][3] ) );
  MXI2X2 U83 ( .A(\u_div/SumTmp[13][2] ), .B(\u_div/PartRem[14][2] ), .S0(
        \u_div/CryTmp[13][6] ), .Y(\u_div/PartRem[13][3] ) );
  MXI2X2 U84 ( .A(\u_div/SumTmp[57][2] ), .B(\u_div/PartRem[58][2] ), .S0(
        \u_div/CryTmp[57][6] ), .Y(\u_div/PartRem[57][3] ) );
  MXI2X2 U85 ( .A(\u_div/SumTmp[15][2] ), .B(\u_div/PartRem[16][2] ), .S0(
        \u_div/CryTmp[15][6] ), .Y(\u_div/PartRem[15][3] ) );
  MXI2X2 U86 ( .A(\u_div/SumTmp[52][2] ), .B(\u_div/PartRem[53][2] ), .S0(
        \u_div/CryTmp[52][6] ), .Y(\u_div/PartRem[52][3] ) );
  MXI2X2 U87 ( .A(\u_div/SumTmp[47][2] ), .B(\u_div/PartRem[48][2] ), .S0(
        \u_div/CryTmp[47][6] ), .Y(\u_div/PartRem[47][3] ) );
  MXI2X2 U88 ( .A(\u_div/SumTmp[42][2] ), .B(\u_div/PartRem[43][2] ), .S0(
        \u_div/CryTmp[42][6] ), .Y(\u_div/PartRem[42][3] ) );
  MXI2X2 U89 ( .A(\u_div/SumTmp[37][2] ), .B(\u_div/PartRem[38][2] ), .S0(
        \u_div/CryTmp[37][6] ), .Y(\u_div/PartRem[37][3] ) );
  MXI2X2 U90 ( .A(\u_div/SumTmp[27][2] ), .B(\u_div/PartRem[28][2] ), .S0(
        \u_div/CryTmp[27][6] ), .Y(\u_div/PartRem[27][3] ) );
  MXI2X2 U91 ( .A(\u_div/SumTmp[22][2] ), .B(\u_div/PartRem[23][2] ), .S0(
        \u_div/CryTmp[22][6] ), .Y(\u_div/PartRem[22][3] ) );
  OR2X2 U92 ( .A(\u_div/PartRem[41][2] ), .B(\u_div/PartRem[41][3] ), .Y(
        \u_div/u_add_PartRem_2_40/n3 ) );
  OR2X2 U93 ( .A(\u_div/PartRem[36][2] ), .B(\u_div/PartRem[36][3] ), .Y(
        \u_div/u_add_PartRem_2_35/n3 ) );
  OR2X2 U94 ( .A(\u_div/PartRem[26][2] ), .B(\u_div/PartRem[26][3] ), .Y(
        \u_div/u_add_PartRem_2_25/n3 ) );
  OR2X2 U95 ( .A(\u_div/PartRem[21][2] ), .B(\u_div/PartRem[21][3] ), .Y(
        \u_div/u_add_PartRem_2_20/n3 ) );
  OR2X2 U96 ( .A(\u_div/PartRem[31][2] ), .B(\u_div/PartRem[31][3] ), .Y(
        \u_div/u_add_PartRem_2_30/n3 ) );
  OR2X2 U97 ( .A(\u_div/PartRem[20][2] ), .B(\u_div/PartRem[20][3] ), .Y(
        \u_div/u_add_PartRem_2_19/n3 ) );
  OR2X2 U98 ( .A(\u_div/PartRem[40][2] ), .B(\u_div/PartRem[40][3] ), .Y(
        \u_div/u_add_PartRem_2_39/n3 ) );
  OR2X2 U99 ( .A(\u_div/PartRem[35][2] ), .B(\u_div/PartRem[35][3] ), .Y(
        \u_div/u_add_PartRem_2_34/n3 ) );
  OR2X2 U100 ( .A(\u_div/PartRem[30][2] ), .B(\u_div/PartRem[30][3] ), .Y(
        \u_div/u_add_PartRem_2_29/n3 ) );
  OR2X2 U101 ( .A(\u_div/PartRem[25][2] ), .B(\u_div/PartRem[25][3] ), .Y(
        \u_div/u_add_PartRem_2_24/n3 ) );
  OR2X2 U102 ( .A(\u_div/PartRem[56][2] ), .B(\u_div/PartRem[56][3] ), .Y(
        \u_div/u_add_PartRem_2_55/n3 ) );
  OR2X2 U103 ( .A(\u_div/PartRem[50][2] ), .B(\u_div/PartRem[50][3] ), .Y(
        \u_div/u_add_PartRem_2_49/n3 ) );
  OR2X2 U104 ( .A(\u_div/PartRem[51][2] ), .B(\u_div/PartRem[51][3] ), .Y(
        \u_div/u_add_PartRem_2_50/n3 ) );
  OR2X2 U105 ( .A(\u_div/PartRem[46][2] ), .B(\u_div/PartRem[46][3] ), .Y(
        \u_div/u_add_PartRem_2_45/n3 ) );
  OR2X2 U106 ( .A(\u_div/PartRem[55][2] ), .B(\u_div/PartRem[55][3] ), .Y(
        \u_div/u_add_PartRem_2_54/n3 ) );
  OR2X2 U107 ( .A(\u_div/PartRem[45][2] ), .B(\u_div/PartRem[45][3] ), .Y(
        \u_div/u_add_PartRem_2_44/n3 ) );
  OR2X2 U108 ( .A(\u_div/PartRem[28][2] ), .B(\u_div/PartRem[28][3] ), .Y(
        \u_div/u_add_PartRem_2_27/n3 ) );
  OR2X2 U109 ( .A(\u_div/PartRem[29][2] ), .B(\u_div/PartRem[29][3] ), .Y(
        \u_div/u_add_PartRem_2_28/n3 ) );
  OR2X2 U110 ( .A(\u_div/PartRem[33][2] ), .B(\u_div/PartRem[33][3] ), .Y(
        \u_div/u_add_PartRem_2_32/n3 ) );
  OR2X2 U111 ( .A(\u_div/PartRem[24][2] ), .B(\u_div/PartRem[24][3] ), .Y(
        \u_div/u_add_PartRem_2_23/n3 ) );
  OR2X2 U112 ( .A(\u_div/PartRem[34][2] ), .B(\u_div/PartRem[34][3] ), .Y(
        \u_div/u_add_PartRem_2_33/n3 ) );
  OR2X2 U113 ( .A(\u_div/PartRem[19][2] ), .B(\u_div/PartRem[19][3] ), .Y(
        \u_div/u_add_PartRem_2_18/n3 ) );
  OR2X2 U114 ( .A(\u_div/PartRem[38][2] ), .B(\u_div/PartRem[38][3] ), .Y(
        \u_div/u_add_PartRem_2_37/n3 ) );
  OR2X2 U115 ( .A(\u_div/PartRem[23][2] ), .B(\u_div/PartRem[23][3] ), .Y(
        \u_div/u_add_PartRem_2_22/n3 ) );
  OR2X2 U116 ( .A(\u_div/PartRem[49][2] ), .B(\u_div/PartRem[49][3] ), .Y(
        \u_div/u_add_PartRem_2_48/n3 ) );
  OR2X2 U117 ( .A(\u_div/PartRem[39][2] ), .B(\u_div/PartRem[39][3] ), .Y(
        \u_div/u_add_PartRem_2_38/n3 ) );
  OR2X2 U118 ( .A(\u_div/PartRem[48][2] ), .B(\u_div/PartRem[48][3] ), .Y(
        \u_div/u_add_PartRem_2_47/n3 ) );
  OR2X2 U119 ( .A(\u_div/PartRem[43][2] ), .B(\u_div/PartRem[43][3] ), .Y(
        \u_div/u_add_PartRem_2_42/n3 ) );
  OR2X2 U120 ( .A(\u_div/PartRem[18][2] ), .B(\u_div/PartRem[18][3] ), .Y(
        \u_div/u_add_PartRem_2_17/n3 ) );
  OR2X2 U121 ( .A(\u_div/PartRem[54][2] ), .B(\u_div/PartRem[54][3] ), .Y(
        \u_div/u_add_PartRem_2_53/n3 ) );
  OR2X2 U122 ( .A(\u_div/PartRem[16][2] ), .B(\u_div/PartRem[16][3] ), .Y(
        \u_div/u_add_PartRem_2_15/n3 ) );
  OR2X2 U123 ( .A(\u_div/PartRem[44][2] ), .B(\u_div/PartRem[44][3] ), .Y(
        \u_div/u_add_PartRem_2_43/n3 ) );
  OR2X2 U124 ( .A(\u_div/PartRem[53][2] ), .B(\u_div/PartRem[53][3] ), .Y(
        \u_div/u_add_PartRem_2_52/n3 ) );
  OR2X2 U125 ( .A(\u_div/PartRem[14][2] ), .B(\u_div/PartRem[14][3] ), .Y(
        \u_div/u_add_PartRem_2_13/n3 ) );
  OR2X2 U126 ( .A(\u_div/PartRem[58][2] ), .B(\u_div/PartRem[58][3] ), .Y(
        \u_div/u_add_PartRem_2_57/n3 ) );
  OR2X2 U127 ( .A(\u_div/PartRem[12][2] ), .B(\u_div/PartRem[12][3] ), .Y(
        \u_div/u_add_PartRem_2_11/n3 ) );
  OR2X2 U128 ( .A(\u_div/PartRem[11][2] ), .B(\u_div/PartRem[11][3] ), .Y(
        \u_div/u_add_PartRem_2_10/n3 ) );
  OR2X2 U129 ( .A(\u_div/PartRem[8][2] ), .B(\u_div/PartRem[8][3] ), .Y(
        \u_div/u_add_PartRem_2_7/n3 ) );
  OR2X2 U130 ( .A(\u_div/PartRem[10][2] ), .B(\u_div/PartRem[10][3] ), .Y(
        \u_div/u_add_PartRem_2_9/n3 ) );
  OR2X2 U131 ( .A(\u_div/PartRem[9][2] ), .B(\u_div/PartRem[9][3] ), .Y(
        \u_div/u_add_PartRem_2_8/n3 ) );
  OR2X2 U132 ( .A(\u_div/PartRem[7][2] ), .B(\u_div/PartRem[7][3] ), .Y(
        \u_div/u_add_PartRem_2_6/n3 ) );
  OR2X2 U133 ( .A(\u_div/PartRem[6][2] ), .B(\u_div/PartRem[6][3] ), .Y(
        \u_div/u_add_PartRem_2_5/n3 ) );
  OR2X2 U134 ( .A(\u_div/PartRem[4][2] ), .B(\u_div/PartRem[4][3] ), .Y(
        \u_div/u_add_PartRem_2_3/n3 ) );
  OR2X2 U135 ( .A(\u_div/PartRem[3][2] ), .B(\u_div/PartRem[3][3] ), .Y(
        \u_div/u_add_PartRem_2_2/n3 ) );
  OR2X2 U136 ( .A(\u_div/PartRem[2][2] ), .B(\u_div/PartRem[2][3] ), .Y(
        \u_div/u_add_PartRem_2_1/n3 ) );
  OR2X2 U137 ( .A(\u_div/PartRem[59][2] ), .B(\u_div/PartRem[59][3] ), .Y(
        \u_div/u_add_PartRem_2_58/n3 ) );
  OR2X1 U138 ( .A(\u_div/PartRem[5][2] ), .B(\u_div/PartRem[5][3] ), .Y(
        \u_div/u_add_PartRem_2_4/n3 ) );
  XNOR2XL U139 ( .A(\u_div/PartRem[64][0] ), .B(n8), .Y(\u_div/SumTmp[59][4] )
         );
  XOR2XL U140 ( .A(\u_div/CryTmp[59][6] ), .B(n3), .Y(\u_div/QInv[59] ) );
  XOR2XL U141 ( .A(\u_div/CryTmp[15][6] ), .B(n4), .Y(\u_div/QInv[15] ) );
  XOR2XL U142 ( .A(\u_div/CryTmp[1][6] ), .B(n4), .Y(\u_div/QInv[1] ) );
  XOR2XL U143 ( .A(\u_div/CryTmp[58][6] ), .B(n5), .Y(\u_div/QInv[58] ) );
  XOR2XL U144 ( .A(\u_div/CryTmp[56][6] ), .B(n3), .Y(\u_div/QInv[56] ) );
  XOR2XL U145 ( .A(\u_div/CryTmp[53][6] ), .B(n3), .Y(\u_div/QInv[53] ) );
  XOR2XL U146 ( .A(\u_div/CryTmp[50][6] ), .B(n3), .Y(\u_div/QInv[50] ) );
  XOR2XL U147 ( .A(\u_div/CryTmp[51][6] ), .B(n4), .Y(\u_div/QInv[51] ) );
  XOR2XL U148 ( .A(\u_div/CryTmp[45][6] ), .B(n3), .Y(\u_div/QInv[45] ) );
  XOR2XL U149 ( .A(\u_div/CryTmp[52][6] ), .B(n5), .Y(\u_div/QInv[52] ) );
  XOR2XL U150 ( .A(\u_div/CryTmp[46][6] ), .B(n4), .Y(\u_div/QInv[46] ) );
  XOR2XL U151 ( .A(\u_div/CryTmp[49][6] ), .B(n4), .Y(\u_div/QInv[49] ) );
  XOR2XL U152 ( .A(\u_div/CryTmp[48][6] ), .B(n3), .Y(\u_div/QInv[48] ) );
  XOR2XL U153 ( .A(\u_div/CryTmp[42][6] ), .B(n3), .Y(\u_div/QInv[42] ) );
  XOR2XL U154 ( .A(\u_div/CryTmp[47][6] ), .B(n5), .Y(\u_div/QInv[47] ) );
  XOR2XL U155 ( .A(\u_div/CryTmp[39][6] ), .B(n5), .Y(\u_div/QInv[39] ) );
  XOR2XL U156 ( .A(\u_div/CryTmp[40][6] ), .B(n4), .Y(\u_div/QInv[40] ) );
  XOR2XL U157 ( .A(\u_div/CryTmp[38][6] ), .B(n4), .Y(\u_div/QInv[38] ) );
  XOR2XL U158 ( .A(\u_div/CryTmp[37][6] ), .B(n3), .Y(\u_div/QInv[37] ) );
  XOR2XL U159 ( .A(\u_div/CryTmp[41][6] ), .B(n5), .Y(\u_div/QInv[41] ) );
  XOR2XL U160 ( .A(\u_div/CryTmp[35][6] ), .B(n4), .Y(\u_div/QInv[35] ) );
  XOR2XL U161 ( .A(\u_div/CryTmp[34][6] ), .B(n5), .Y(\u_div/QInv[34] ) );
  XOR2XL U162 ( .A(\u_div/CryTmp[33][6] ), .B(n4), .Y(\u_div/QInv[33] ) );
  XOR2XL U163 ( .A(\u_div/CryTmp[36][6] ), .B(n5), .Y(\u_div/QInv[36] ) );
  XOR2XL U164 ( .A(\u_div/CryTmp[30][6] ), .B(n4), .Y(\u_div/QInv[30] ) );
  XOR2XL U165 ( .A(\u_div/CryTmp[28][6] ), .B(n4), .Y(\u_div/QInv[28] ) );
  XOR2XL U166 ( .A(\u_div/CryTmp[29][6] ), .B(n5), .Y(\u_div/QInv[29] ) );
  XOR2XL U167 ( .A(\u_div/CryTmp[27][6] ), .B(n3), .Y(\u_div/QInv[27] ) );
  XOR2XL U168 ( .A(\u_div/CryTmp[25][6] ), .B(n4), .Y(\u_div/QInv[25] ) );
  XOR2XL U169 ( .A(\u_div/CryTmp[26][6] ), .B(n5), .Y(\u_div/QInv[26] ) );
  XOR2XL U170 ( .A(\u_div/CryTmp[24][6] ), .B(n3), .Y(\u_div/QInv[24] ) );
  XOR2XL U171 ( .A(\u_div/CryTmp[22][6] ), .B(n4), .Y(\u_div/QInv[22] ) );
  XOR2XL U172 ( .A(\u_div/CryTmp[21][6] ), .B(n3), .Y(\u_div/QInv[21] ) );
  XOR2XL U173 ( .A(\u_div/CryTmp[23][6] ), .B(n5), .Y(\u_div/QInv[23] ) );
  XOR2XL U174 ( .A(\u_div/CryTmp[20][6] ), .B(n5), .Y(\u_div/QInv[20] ) );
  XOR2XL U175 ( .A(\u_div/CryTmp[19][6] ), .B(n3), .Y(\u_div/QInv[19] ) );
  XOR2XL U176 ( .A(\u_div/CryTmp[10][6] ), .B(n5), .Y(\u_div/QInv[10] ) );
  XOR2XL U177 ( .A(\u_div/CryTmp[16][6] ), .B(n5), .Y(\u_div/QInv[16] ) );
  INVXL U178 ( .A(\u_div/PartRem[59][2] ), .Y(\u_div/SumTmp[58][2] ) );
  INVXL U179 ( .A(\u_div/PartRem[54][2] ), .Y(\u_div/SumTmp[53][2] ) );
  INVXL U180 ( .A(\u_div/PartRem[49][2] ), .Y(\u_div/SumTmp[48][2] ) );
  INVXL U181 ( .A(\u_div/PartRem[44][2] ), .Y(\u_div/SumTmp[43][2] ) );
  INVXL U182 ( .A(\u_div/PartRem[39][2] ), .Y(\u_div/SumTmp[38][2] ) );
  INVXL U183 ( .A(\u_div/PartRem[34][2] ), .Y(\u_div/SumTmp[33][2] ) );
  INVXL U184 ( .A(\u_div/PartRem[29][2] ), .Y(\u_div/SumTmp[28][2] ) );
  INVXL U185 ( .A(\u_div/PartRem[24][2] ), .Y(\u_div/SumTmp[23][2] ) );
  INVXL U186 ( .A(\u_div/PartRem[19][2] ), .Y(\u_div/SumTmp[18][2] ) );
  INVX3 U187 ( .A(n2), .Y(n3) );
  MXI2X1 U188 ( .A(\u_div/SumTmp[1][1] ), .B(\u_div/SumTmp[1][1] ), .S0(
        \u_div/CryTmp[1][6] ), .Y(n1) );
  CLKINVX1 U189 ( .A(\u_div/QInv[63] ), .Y(n2) );
  MXI2X1 U190 ( .A(\u_div/SumTmp[2][2] ), .B(\u_div/PartRem[3][2] ), .S0(
        \u_div/CryTmp[2][6] ), .Y(\u_div/PartRem[2][3] ) );
  CLKINVX1 U191 ( .A(\u_div/PartRem[3][2] ), .Y(\u_div/SumTmp[2][2] ) );
  MXI2X1 U192 ( .A(\u_div/SumTmp[58][2] ), .B(\u_div/PartRem[59][2] ), .S0(
        \u_div/CryTmp[58][6] ), .Y(\u_div/PartRem[58][3] ) );
  CLKINVX1 U193 ( .A(\u_div/PartRem[58][2] ), .Y(\u_div/SumTmp[57][2] ) );
  MXI2X1 U194 ( .A(\u_div/SumTmp[56][2] ), .B(\u_div/PartRem[57][2] ), .S0(
        \u_div/CryTmp[56][6] ), .Y(\u_div/PartRem[56][3] ) );
  CLKINVX1 U195 ( .A(\u_div/PartRem[57][2] ), .Y(\u_div/SumTmp[56][2] ) );
  MXI2X1 U196 ( .A(\u_div/SumTmp[55][2] ), .B(\u_div/PartRem[56][2] ), .S0(
        \u_div/CryTmp[55][6] ), .Y(\u_div/PartRem[55][3] ) );
  CLKINVX1 U197 ( .A(\u_div/PartRem[56][2] ), .Y(\u_div/SumTmp[55][2] ) );
  MXI2X1 U198 ( .A(\u_div/SumTmp[53][2] ), .B(\u_div/PartRem[54][2] ), .S0(
        \u_div/CryTmp[53][6] ), .Y(\u_div/PartRem[53][3] ) );
  CLKINVX1 U199 ( .A(\u_div/PartRem[53][2] ), .Y(\u_div/SumTmp[52][2] ) );
  MXI2X1 U200 ( .A(\u_div/SumTmp[51][2] ), .B(\u_div/PartRem[52][2] ), .S0(
        \u_div/CryTmp[51][6] ), .Y(\u_div/PartRem[51][3] ) );
  CLKINVX1 U201 ( .A(\u_div/PartRem[52][2] ), .Y(\u_div/SumTmp[51][2] ) );
  MXI2X1 U202 ( .A(\u_div/SumTmp[50][2] ), .B(\u_div/PartRem[51][2] ), .S0(
        \u_div/CryTmp[50][6] ), .Y(\u_div/PartRem[50][3] ) );
  CLKINVX1 U203 ( .A(\u_div/PartRem[51][2] ), .Y(\u_div/SumTmp[50][2] ) );
  MXI2X1 U204 ( .A(\u_div/SumTmp[48][2] ), .B(\u_div/PartRem[49][2] ), .S0(
        \u_div/CryTmp[48][6] ), .Y(\u_div/PartRem[48][3] ) );
  CLKINVX1 U205 ( .A(\u_div/PartRem[48][2] ), .Y(\u_div/SumTmp[47][2] ) );
  MXI2X1 U206 ( .A(\u_div/SumTmp[46][2] ), .B(\u_div/PartRem[47][2] ), .S0(
        \u_div/CryTmp[46][6] ), .Y(\u_div/PartRem[46][3] ) );
  CLKINVX1 U207 ( .A(\u_div/PartRem[47][2] ), .Y(\u_div/SumTmp[46][2] ) );
  MXI2X1 U208 ( .A(\u_div/SumTmp[45][2] ), .B(\u_div/PartRem[46][2] ), .S0(
        \u_div/CryTmp[45][6] ), .Y(\u_div/PartRem[45][3] ) );
  CLKINVX1 U209 ( .A(\u_div/PartRem[46][2] ), .Y(\u_div/SumTmp[45][2] ) );
  MXI2X1 U210 ( .A(\u_div/SumTmp[43][2] ), .B(\u_div/PartRem[44][2] ), .S0(
        \u_div/CryTmp[43][6] ), .Y(\u_div/PartRem[43][3] ) );
  CLKINVX1 U211 ( .A(\u_div/PartRem[43][2] ), .Y(\u_div/SumTmp[42][2] ) );
  MXI2X1 U212 ( .A(\u_div/SumTmp[41][2] ), .B(\u_div/PartRem[42][2] ), .S0(
        \u_div/CryTmp[41][6] ), .Y(\u_div/PartRem[41][3] ) );
  CLKINVX1 U213 ( .A(\u_div/PartRem[42][2] ), .Y(\u_div/SumTmp[41][2] ) );
  MXI2X1 U214 ( .A(\u_div/SumTmp[40][2] ), .B(\u_div/PartRem[41][2] ), .S0(
        \u_div/CryTmp[40][6] ), .Y(\u_div/PartRem[40][3] ) );
  CLKINVX1 U215 ( .A(\u_div/PartRem[41][2] ), .Y(\u_div/SumTmp[40][2] ) );
  MXI2X1 U216 ( .A(\u_div/SumTmp[38][2] ), .B(\u_div/PartRem[39][2] ), .S0(
        \u_div/CryTmp[38][6] ), .Y(\u_div/PartRem[38][3] ) );
  CLKINVX1 U217 ( .A(\u_div/PartRem[38][2] ), .Y(\u_div/SumTmp[37][2] ) );
  MXI2X1 U218 ( .A(\u_div/SumTmp[36][2] ), .B(\u_div/PartRem[37][2] ), .S0(
        \u_div/CryTmp[36][6] ), .Y(\u_div/PartRem[36][3] ) );
  CLKINVX1 U219 ( .A(\u_div/PartRem[37][2] ), .Y(\u_div/SumTmp[36][2] ) );
  MXI2X1 U220 ( .A(\u_div/SumTmp[35][2] ), .B(\u_div/PartRem[36][2] ), .S0(
        \u_div/CryTmp[35][6] ), .Y(\u_div/PartRem[35][3] ) );
  CLKINVX1 U221 ( .A(\u_div/PartRem[36][2] ), .Y(\u_div/SumTmp[35][2] ) );
  MXI2X1 U222 ( .A(\u_div/SumTmp[33][2] ), .B(\u_div/PartRem[34][2] ), .S0(
        \u_div/CryTmp[33][6] ), .Y(\u_div/PartRem[33][3] ) );
  CLKINVX1 U223 ( .A(\u_div/PartRem[33][2] ), .Y(\u_div/SumTmp[32][2] ) );
  MXI2X1 U224 ( .A(\u_div/SumTmp[31][2] ), .B(\u_div/PartRem[32][2] ), .S0(
        \u_div/CryTmp[31][6] ), .Y(\u_div/PartRem[31][3] ) );
  CLKINVX1 U225 ( .A(\u_div/PartRem[32][2] ), .Y(\u_div/SumTmp[31][2] ) );
  MXI2X1 U226 ( .A(\u_div/SumTmp[30][2] ), .B(\u_div/PartRem[31][2] ), .S0(
        \u_div/CryTmp[30][6] ), .Y(\u_div/PartRem[30][3] ) );
  CLKINVX1 U227 ( .A(\u_div/PartRem[31][2] ), .Y(\u_div/SumTmp[30][2] ) );
  MXI2X1 U228 ( .A(\u_div/SumTmp[28][2] ), .B(\u_div/PartRem[29][2] ), .S0(
        \u_div/CryTmp[28][6] ), .Y(\u_div/PartRem[28][3] ) );
  CLKINVX1 U229 ( .A(\u_div/PartRem[28][2] ), .Y(\u_div/SumTmp[27][2] ) );
  MXI2X1 U230 ( .A(\u_div/SumTmp[26][2] ), .B(\u_div/PartRem[27][2] ), .S0(
        \u_div/CryTmp[26][6] ), .Y(\u_div/PartRem[26][3] ) );
  CLKINVX1 U231 ( .A(\u_div/PartRem[27][2] ), .Y(\u_div/SumTmp[26][2] ) );
  MXI2X1 U232 ( .A(\u_div/SumTmp[25][2] ), .B(\u_div/PartRem[26][2] ), .S0(
        \u_div/CryTmp[25][6] ), .Y(\u_div/PartRem[25][3] ) );
  CLKINVX1 U233 ( .A(\u_div/PartRem[26][2] ), .Y(\u_div/SumTmp[25][2] ) );
  MXI2X1 U234 ( .A(\u_div/SumTmp[23][2] ), .B(\u_div/PartRem[24][2] ), .S0(
        \u_div/CryTmp[23][6] ), .Y(\u_div/PartRem[23][3] ) );
  CLKINVX1 U235 ( .A(\u_div/PartRem[23][2] ), .Y(\u_div/SumTmp[22][2] ) );
  MXI2X1 U236 ( .A(\u_div/SumTmp[21][2] ), .B(\u_div/PartRem[22][2] ), .S0(
        \u_div/CryTmp[21][6] ), .Y(\u_div/PartRem[21][3] ) );
  CLKINVX1 U237 ( .A(\u_div/PartRem[22][2] ), .Y(\u_div/SumTmp[21][2] ) );
  MXI2X1 U238 ( .A(\u_div/SumTmp[20][2] ), .B(\u_div/PartRem[21][2] ), .S0(
        \u_div/CryTmp[20][6] ), .Y(\u_div/PartRem[20][3] ) );
  CLKINVX1 U239 ( .A(\u_div/PartRem[21][2] ), .Y(\u_div/SumTmp[20][2] ) );
  MXI2X1 U240 ( .A(\u_div/SumTmp[18][2] ), .B(\u_div/PartRem[19][2] ), .S0(
        \u_div/CryTmp[18][6] ), .Y(\u_div/PartRem[18][3] ) );
  CLKINVX1 U241 ( .A(\u_div/PartRem[18][2] ), .Y(\u_div/SumTmp[17][2] ) );
  MXI2X1 U242 ( .A(\u_div/SumTmp[16][2] ), .B(\u_div/PartRem[17][2] ), .S0(
        \u_div/CryTmp[16][6] ), .Y(\u_div/PartRem[16][3] ) );
  CLKINVX1 U243 ( .A(\u_div/PartRem[17][2] ), .Y(\u_div/SumTmp[16][2] ) );
  MXI2X1 U244 ( .A(\u_div/SumTmp[14][2] ), .B(\u_div/PartRem[15][2] ), .S0(
        \u_div/CryTmp[14][6] ), .Y(\u_div/PartRem[14][3] ) );
  CLKINVX1 U245 ( .A(\u_div/PartRem[15][2] ), .Y(\u_div/SumTmp[14][2] ) );
  MXI2X1 U246 ( .A(\u_div/SumTmp[11][2] ), .B(\u_div/PartRem[12][2] ), .S0(
        \u_div/CryTmp[11][6] ), .Y(\u_div/PartRem[11][3] ) );
  CLKINVX1 U247 ( .A(\u_div/PartRem[12][2] ), .Y(\u_div/SumTmp[11][2] ) );
  MXI2X1 U248 ( .A(\u_div/SumTmp[6][2] ), .B(\u_div/PartRem[7][2] ), .S0(
        \u_div/CryTmp[6][6] ), .Y(\u_div/PartRem[6][3] ) );
  CLKINVX1 U249 ( .A(\u_div/PartRem[7][2] ), .Y(\u_div/SumTmp[6][2] ) );
  MXI2X1 U250 ( .A(\u_div/SumTmp[10][2] ), .B(\u_div/PartRem[11][2] ), .S0(
        \u_div/CryTmp[10][6] ), .Y(\u_div/PartRem[10][3] ) );
  CLKINVX1 U251 ( .A(\u_div/PartRem[11][2] ), .Y(\u_div/SumTmp[10][2] ) );
  MXI2X1 U252 ( .A(\u_div/SumTmp[5][2] ), .B(\u_div/PartRem[6][2] ), .S0(
        \u_div/CryTmp[5][6] ), .Y(\u_div/PartRem[5][3] ) );
  CLKINVX1 U253 ( .A(\u_div/PartRem[6][2] ), .Y(\u_div/SumTmp[5][2] ) );
  CLKINVX1 U254 ( .A(\u_div/PartRem[16][2] ), .Y(\u_div/SumTmp[15][2] ) );
  CLKINVX1 U255 ( .A(\u_div/PartRem[14][2] ), .Y(\u_div/SumTmp[13][2] ) );
  MXI2X1 U256 ( .A(\u_div/SumTmp[12][2] ), .B(\u_div/PartRem[13][2] ), .S0(
        \u_div/CryTmp[12][6] ), .Y(\u_div/PartRem[12][3] ) );
  CLKINVX1 U257 ( .A(\u_div/PartRem[13][2] ), .Y(\u_div/SumTmp[12][2] ) );
  MXI2X1 U258 ( .A(\u_div/SumTmp[9][2] ), .B(\u_div/PartRem[10][2] ), .S0(
        \u_div/CryTmp[9][6] ), .Y(\u_div/PartRem[9][3] ) );
  CLKINVX1 U259 ( .A(\u_div/PartRem[10][2] ), .Y(\u_div/SumTmp[9][2] ) );
  MXI2X1 U260 ( .A(\u_div/SumTmp[8][2] ), .B(\u_div/PartRem[9][2] ), .S0(
        \u_div/CryTmp[8][6] ), .Y(\u_div/PartRem[8][3] ) );
  CLKINVX1 U261 ( .A(\u_div/PartRem[9][2] ), .Y(\u_div/SumTmp[8][2] ) );
  MXI2X1 U262 ( .A(\u_div/SumTmp[7][2] ), .B(\u_div/PartRem[8][2] ), .S0(
        \u_div/CryTmp[7][6] ), .Y(\u_div/PartRem[7][3] ) );
  CLKINVX1 U263 ( .A(\u_div/PartRem[8][2] ), .Y(\u_div/SumTmp[7][2] ) );
  MXI2X1 U264 ( .A(\u_div/SumTmp[4][2] ), .B(\u_div/PartRem[5][2] ), .S0(
        \u_div/CryTmp[4][6] ), .Y(\u_div/PartRem[4][3] ) );
  CLKINVX1 U265 ( .A(\u_div/PartRem[5][2] ), .Y(\u_div/SumTmp[4][2] ) );
  MXI2X1 U266 ( .A(\u_div/SumTmp[3][2] ), .B(\u_div/PartRem[4][2] ), .S0(
        \u_div/CryTmp[3][6] ), .Y(\u_div/PartRem[3][3] ) );
  CLKINVX1 U267 ( .A(\u_div/PartRem[4][2] ), .Y(\u_div/SumTmp[3][2] ) );
  MXI2X1 U268 ( .A(n7), .B(\u_div/PartRem[62][0] ), .S0(\u_div/CryTmp[59][6] ), 
        .Y(\u_div/PartRem[59][3] ) );
  CLKINVX1 U269 ( .A(\u_div/PartRem[62][0] ), .Y(n7) );
  MXI2X1 U270 ( .A(\u_div/SumTmp[54][2] ), .B(\u_div/PartRem[55][2] ), .S0(
        \u_div/CryTmp[54][6] ), .Y(\u_div/PartRem[54][3] ) );
  CLKINVX1 U271 ( .A(\u_div/PartRem[55][2] ), .Y(\u_div/SumTmp[54][2] ) );
  MXI2X1 U272 ( .A(\u_div/SumTmp[49][2] ), .B(\u_div/PartRem[50][2] ), .S0(
        \u_div/CryTmp[49][6] ), .Y(\u_div/PartRem[49][3] ) );
  CLKINVX1 U273 ( .A(\u_div/PartRem[50][2] ), .Y(\u_div/SumTmp[49][2] ) );
  MXI2X1 U274 ( .A(\u_div/SumTmp[44][2] ), .B(\u_div/PartRem[45][2] ), .S0(
        \u_div/CryTmp[44][6] ), .Y(\u_div/PartRem[44][3] ) );
  CLKINVX1 U275 ( .A(\u_div/PartRem[45][2] ), .Y(\u_div/SumTmp[44][2] ) );
  MXI2X1 U276 ( .A(\u_div/SumTmp[39][2] ), .B(\u_div/PartRem[40][2] ), .S0(
        \u_div/CryTmp[39][6] ), .Y(\u_div/PartRem[39][3] ) );
  CLKINVX1 U277 ( .A(\u_div/PartRem[40][2] ), .Y(\u_div/SumTmp[39][2] ) );
  MXI2X1 U278 ( .A(\u_div/SumTmp[34][2] ), .B(\u_div/PartRem[35][2] ), .S0(
        \u_div/CryTmp[34][6] ), .Y(\u_div/PartRem[34][3] ) );
  CLKINVX1 U279 ( .A(\u_div/PartRem[35][2] ), .Y(\u_div/SumTmp[34][2] ) );
  MXI2X1 U280 ( .A(\u_div/SumTmp[29][2] ), .B(\u_div/PartRem[30][2] ), .S0(
        \u_div/CryTmp[29][6] ), .Y(\u_div/PartRem[29][3] ) );
  CLKINVX1 U281 ( .A(\u_div/PartRem[30][2] ), .Y(\u_div/SumTmp[29][2] ) );
  MXI2X1 U282 ( .A(\u_div/SumTmp[24][2] ), .B(\u_div/PartRem[25][2] ), .S0(
        \u_div/CryTmp[24][6] ), .Y(\u_div/PartRem[24][3] ) );
  CLKINVX1 U283 ( .A(\u_div/PartRem[25][2] ), .Y(\u_div/SumTmp[24][2] ) );
  MXI2X1 U284 ( .A(\u_div/SumTmp[19][2] ), .B(\u_div/PartRem[20][2] ), .S0(
        \u_div/CryTmp[19][6] ), .Y(\u_div/PartRem[19][3] ) );
  CLKINVX1 U285 ( .A(\u_div/PartRem[20][2] ), .Y(\u_div/SumTmp[19][2] ) );
  CLKINVX1 U286 ( .A(\u_div/PartRem[2][2] ), .Y(\u_div/SumTmp[1][2] ) );
  INVX4 U287 ( .A(n2), .Y(n4) );
  INVX4 U288 ( .A(n2), .Y(n5) );
  XOR2XL U289 ( .A(\u_div/CryTmp[14][6] ), .B(n5), .Y(\u_div/QInv[14] ) );
  XOR2XL U290 ( .A(\u_div/CryTmp[12][6] ), .B(n5), .Y(\u_div/QInv[12] ) );
  XOR2XL U291 ( .A(\u_div/CryTmp[11][6] ), .B(n4), .Y(\u_div/QInv[11] ) );
  XOR2XL U292 ( .A(\u_div/CryTmp[9][6] ), .B(n3), .Y(\u_div/QInv[9] ) );
  XOR2XL U293 ( .A(\u_div/CryTmp[8][6] ), .B(n3), .Y(\u_div/QInv[8] ) );
  XOR2XL U294 ( .A(\u_div/CryTmp[7][6] ), .B(n4), .Y(\u_div/QInv[7] ) );
  XOR2XL U295 ( .A(\u_div/CryTmp[6][6] ), .B(n5), .Y(\u_div/QInv[6] ) );
  XOR2XL U296 ( .A(\u_div/CryTmp[4][6] ), .B(n5), .Y(\u_div/QInv[4] ) );
  XOR2XL U297 ( .A(\u_div/CryTmp[3][6] ), .B(n3), .Y(\u_div/QInv[3] ) );
  XOR2XL U298 ( .A(\u_div/CryTmp[2][6] ), .B(n3), .Y(\u_div/QInv[2] ) );
  XNOR2X1 U299 ( .A(\u_div/PartRem[59][3] ), .B(\u_div/PartRem[59][2] ), .Y(
        \u_div/SumTmp[58][3] ) );
  XNOR2X1 U300 ( .A(\u_div/PartRem[58][3] ), .B(\u_div/PartRem[58][2] ), .Y(
        \u_div/SumTmp[57][3] ) );
  OR2X1 U301 ( .A(\u_div/PartRem[57][5] ), .B(\u_div/u_add_PartRem_2_56/n2 ), 
        .Y(\u_div/CryTmp[56][6] ) );
  XNOR2X1 U302 ( .A(\u_div/PartRem[57][3] ), .B(\u_div/PartRem[57][2] ), .Y(
        \u_div/SumTmp[56][3] ) );
  OR2X1 U303 ( .A(\u_div/PartRem[57][2] ), .B(\u_div/PartRem[57][3] ), .Y(
        \u_div/u_add_PartRem_2_56/n3 ) );
  OR2X1 U304 ( .A(\u_div/PartRem[56][5] ), .B(\u_div/u_add_PartRem_2_55/n2 ), 
        .Y(\u_div/CryTmp[55][6] ) );
  XNOR2X1 U305 ( .A(\u_div/PartRem[56][3] ), .B(\u_div/PartRem[56][2] ), .Y(
        \u_div/SumTmp[55][3] ) );
  XNOR2X1 U306 ( .A(\u_div/PartRem[55][3] ), .B(\u_div/PartRem[55][2] ), .Y(
        \u_div/SumTmp[54][3] ) );
  OR2X1 U307 ( .A(\u_div/PartRem[54][5] ), .B(\u_div/u_add_PartRem_2_53/n2 ), 
        .Y(\u_div/CryTmp[53][6] ) );
  XNOR2X1 U308 ( .A(\u_div/PartRem[54][3] ), .B(\u_div/PartRem[54][2] ), .Y(
        \u_div/SumTmp[53][3] ) );
  OR2X1 U309 ( .A(\u_div/PartRem[53][5] ), .B(\u_div/u_add_PartRem_2_52/n2 ), 
        .Y(\u_div/CryTmp[52][6] ) );
  XNOR2X1 U310 ( .A(\u_div/PartRem[53][3] ), .B(\u_div/PartRem[53][2] ), .Y(
        \u_div/SumTmp[52][3] ) );
  OR2X1 U311 ( .A(\u_div/PartRem[52][5] ), .B(\u_div/u_add_PartRem_2_51/n2 ), 
        .Y(\u_div/CryTmp[51][6] ) );
  XNOR2X1 U312 ( .A(\u_div/PartRem[52][3] ), .B(\u_div/PartRem[52][2] ), .Y(
        \u_div/SumTmp[51][3] ) );
  OR2X1 U313 ( .A(\u_div/PartRem[52][2] ), .B(\u_div/PartRem[52][3] ), .Y(
        \u_div/u_add_PartRem_2_51/n3 ) );
  OR2X1 U314 ( .A(\u_div/PartRem[51][5] ), .B(\u_div/u_add_PartRem_2_50/n2 ), 
        .Y(\u_div/CryTmp[50][6] ) );
  XNOR2X1 U315 ( .A(\u_div/PartRem[51][3] ), .B(\u_div/PartRem[51][2] ), .Y(
        \u_div/SumTmp[50][3] ) );
  XNOR2X1 U316 ( .A(\u_div/PartRem[50][3] ), .B(\u_div/PartRem[50][2] ), .Y(
        \u_div/SumTmp[49][3] ) );
  OR2X1 U317 ( .A(\u_div/PartRem[49][5] ), .B(\u_div/u_add_PartRem_2_48/n2 ), 
        .Y(\u_div/CryTmp[48][6] ) );
  XNOR2X1 U318 ( .A(\u_div/PartRem[49][3] ), .B(\u_div/PartRem[49][2] ), .Y(
        \u_div/SumTmp[48][3] ) );
  XNOR2X1 U319 ( .A(\u_div/PartRem[48][3] ), .B(\u_div/PartRem[48][2] ), .Y(
        \u_div/SumTmp[47][3] ) );
  OR2X1 U320 ( .A(\u_div/PartRem[47][5] ), .B(\u_div/u_add_PartRem_2_46/n2 ), 
        .Y(\u_div/CryTmp[46][6] ) );
  XNOR2X1 U321 ( .A(\u_div/PartRem[47][3] ), .B(\u_div/PartRem[47][2] ), .Y(
        \u_div/SumTmp[46][3] ) );
  OR2X1 U322 ( .A(\u_div/PartRem[47][2] ), .B(\u_div/PartRem[47][3] ), .Y(
        \u_div/u_add_PartRem_2_46/n3 ) );
  OR2X1 U323 ( .A(\u_div/PartRem[46][5] ), .B(\u_div/u_add_PartRem_2_45/n2 ), 
        .Y(\u_div/CryTmp[45][6] ) );
  XNOR2X1 U324 ( .A(\u_div/PartRem[46][3] ), .B(\u_div/PartRem[46][2] ), .Y(
        \u_div/SumTmp[45][3] ) );
  XNOR2X1 U325 ( .A(\u_div/PartRem[45][3] ), .B(\u_div/PartRem[45][2] ), .Y(
        \u_div/SumTmp[44][3] ) );
  OR2X1 U326 ( .A(\u_div/PartRem[44][5] ), .B(\u_div/u_add_PartRem_2_43/n2 ), 
        .Y(\u_div/CryTmp[43][6] ) );
  XNOR2X1 U327 ( .A(\u_div/PartRem[44][3] ), .B(\u_div/PartRem[44][2] ), .Y(
        \u_div/SumTmp[43][3] ) );
  XNOR2X1 U328 ( .A(\u_div/PartRem[43][3] ), .B(\u_div/PartRem[43][2] ), .Y(
        \u_div/SumTmp[42][3] ) );
  OR2X1 U329 ( .A(\u_div/PartRem[42][5] ), .B(\u_div/u_add_PartRem_2_41/n2 ), 
        .Y(\u_div/CryTmp[41][6] ) );
  XNOR2X1 U330 ( .A(\u_div/PartRem[42][3] ), .B(\u_div/PartRem[42][2] ), .Y(
        \u_div/SumTmp[41][3] ) );
  OR2X1 U331 ( .A(\u_div/PartRem[42][2] ), .B(\u_div/PartRem[42][3] ), .Y(
        \u_div/u_add_PartRem_2_41/n3 ) );
  OR2X1 U332 ( .A(\u_div/PartRem[41][5] ), .B(\u_div/u_add_PartRem_2_40/n2 ), 
        .Y(\u_div/CryTmp[40][6] ) );
  XNOR2X1 U333 ( .A(\u_div/PartRem[41][3] ), .B(\u_div/PartRem[41][2] ), .Y(
        \u_div/SumTmp[40][3] ) );
  XNOR2X1 U334 ( .A(\u_div/PartRem[40][3] ), .B(\u_div/PartRem[40][2] ), .Y(
        \u_div/SumTmp[39][3] ) );
  OR2X1 U335 ( .A(\u_div/PartRem[39][5] ), .B(\u_div/u_add_PartRem_2_38/n2 ), 
        .Y(\u_div/CryTmp[38][6] ) );
  XNOR2X1 U336 ( .A(\u_div/PartRem[39][3] ), .B(\u_div/PartRem[39][2] ), .Y(
        \u_div/SumTmp[38][3] ) );
  XNOR2X1 U337 ( .A(\u_div/PartRem[38][3] ), .B(\u_div/PartRem[38][2] ), .Y(
        \u_div/SumTmp[37][3] ) );
  OR2X1 U338 ( .A(\u_div/PartRem[37][5] ), .B(\u_div/u_add_PartRem_2_36/n2 ), 
        .Y(\u_div/CryTmp[36][6] ) );
  XNOR2X1 U339 ( .A(\u_div/PartRem[37][3] ), .B(\u_div/PartRem[37][2] ), .Y(
        \u_div/SumTmp[36][3] ) );
  OR2X1 U340 ( .A(\u_div/PartRem[37][2] ), .B(\u_div/PartRem[37][3] ), .Y(
        \u_div/u_add_PartRem_2_36/n3 ) );
  OR2X1 U341 ( .A(\u_div/PartRem[36][5] ), .B(\u_div/u_add_PartRem_2_35/n2 ), 
        .Y(\u_div/CryTmp[35][6] ) );
  XNOR2X1 U342 ( .A(\u_div/PartRem[36][3] ), .B(\u_div/PartRem[36][2] ), .Y(
        \u_div/SumTmp[35][3] ) );
  XNOR2X1 U343 ( .A(\u_div/PartRem[35][3] ), .B(\u_div/PartRem[35][2] ), .Y(
        \u_div/SumTmp[34][3] ) );
  OR2X1 U344 ( .A(\u_div/PartRem[34][5] ), .B(\u_div/u_add_PartRem_2_33/n2 ), 
        .Y(\u_div/CryTmp[33][6] ) );
  XNOR2X1 U345 ( .A(\u_div/PartRem[34][3] ), .B(\u_div/PartRem[34][2] ), .Y(
        \u_div/SumTmp[33][3] ) );
  XNOR2X1 U346 ( .A(\u_div/PartRem[33][3] ), .B(\u_div/PartRem[33][2] ), .Y(
        \u_div/SumTmp[32][3] ) );
  OR2X1 U347 ( .A(\u_div/PartRem[32][5] ), .B(\u_div/u_add_PartRem_2_31/n2 ), 
        .Y(\u_div/CryTmp[31][6] ) );
  XNOR2X1 U348 ( .A(\u_div/PartRem[32][3] ), .B(\u_div/PartRem[32][2] ), .Y(
        \u_div/SumTmp[31][3] ) );
  OR2X1 U349 ( .A(\u_div/PartRem[32][2] ), .B(\u_div/PartRem[32][3] ), .Y(
        \u_div/u_add_PartRem_2_31/n3 ) );
  OR2X1 U350 ( .A(\u_div/PartRem[31][5] ), .B(\u_div/u_add_PartRem_2_30/n2 ), 
        .Y(\u_div/CryTmp[30][6] ) );
  XNOR2X1 U351 ( .A(\u_div/PartRem[31][3] ), .B(\u_div/PartRem[31][2] ), .Y(
        \u_div/SumTmp[30][3] ) );
  XNOR2X1 U352 ( .A(\u_div/PartRem[30][3] ), .B(\u_div/PartRem[30][2] ), .Y(
        \u_div/SumTmp[29][3] ) );
  OR2X1 U353 ( .A(\u_div/PartRem[29][5] ), .B(\u_div/u_add_PartRem_2_28/n2 ), 
        .Y(\u_div/CryTmp[28][6] ) );
  XNOR2X1 U354 ( .A(\u_div/PartRem[29][3] ), .B(\u_div/PartRem[29][2] ), .Y(
        \u_div/SumTmp[28][3] ) );
  XNOR2X1 U355 ( .A(\u_div/PartRem[28][3] ), .B(\u_div/PartRem[28][2] ), .Y(
        \u_div/SumTmp[27][3] ) );
  OR2X1 U356 ( .A(\u_div/PartRem[27][5] ), .B(\u_div/u_add_PartRem_2_26/n2 ), 
        .Y(\u_div/CryTmp[26][6] ) );
  XNOR2X1 U357 ( .A(\u_div/PartRem[27][3] ), .B(\u_div/PartRem[27][2] ), .Y(
        \u_div/SumTmp[26][3] ) );
  OR2X1 U358 ( .A(\u_div/PartRem[27][2] ), .B(\u_div/PartRem[27][3] ), .Y(
        \u_div/u_add_PartRem_2_26/n3 ) );
  OR2X1 U359 ( .A(\u_div/PartRem[26][5] ), .B(\u_div/u_add_PartRem_2_25/n2 ), 
        .Y(\u_div/CryTmp[25][6] ) );
  XNOR2X1 U360 ( .A(\u_div/PartRem[26][3] ), .B(\u_div/PartRem[26][2] ), .Y(
        \u_div/SumTmp[25][3] ) );
  XNOR2X1 U361 ( .A(\u_div/PartRem[25][3] ), .B(\u_div/PartRem[25][2] ), .Y(
        \u_div/SumTmp[24][3] ) );
  OR2X1 U362 ( .A(\u_div/PartRem[24][5] ), .B(\u_div/u_add_PartRem_2_23/n2 ), 
        .Y(\u_div/CryTmp[23][6] ) );
  XNOR2X1 U363 ( .A(\u_div/PartRem[24][3] ), .B(\u_div/PartRem[24][2] ), .Y(
        \u_div/SumTmp[23][3] ) );
  XNOR2X1 U364 ( .A(\u_div/PartRem[23][3] ), .B(\u_div/PartRem[23][2] ), .Y(
        \u_div/SumTmp[22][3] ) );
  OR2X1 U365 ( .A(\u_div/PartRem[22][5] ), .B(\u_div/u_add_PartRem_2_21/n2 ), 
        .Y(\u_div/CryTmp[21][6] ) );
  XNOR2X1 U366 ( .A(\u_div/PartRem[22][3] ), .B(\u_div/PartRem[22][2] ), .Y(
        \u_div/SumTmp[21][3] ) );
  OR2X1 U367 ( .A(\u_div/PartRem[22][2] ), .B(\u_div/PartRem[22][3] ), .Y(
        \u_div/u_add_PartRem_2_21/n3 ) );
  OR2X1 U368 ( .A(\u_div/PartRem[21][5] ), .B(\u_div/u_add_PartRem_2_20/n2 ), 
        .Y(\u_div/CryTmp[20][6] ) );
  XNOR2X1 U369 ( .A(\u_div/PartRem[21][3] ), .B(\u_div/PartRem[21][2] ), .Y(
        \u_div/SumTmp[20][3] ) );
  XNOR2X1 U370 ( .A(\u_div/PartRem[20][3] ), .B(\u_div/PartRem[20][2] ), .Y(
        \u_div/SumTmp[19][3] ) );
  OR2X1 U371 ( .A(\u_div/PartRem[19][5] ), .B(\u_div/u_add_PartRem_2_18/n2 ), 
        .Y(\u_div/CryTmp[18][6] ) );
  XNOR2X1 U372 ( .A(\u_div/PartRem[19][3] ), .B(\u_div/PartRem[19][2] ), .Y(
        \u_div/SumTmp[18][3] ) );
  XNOR2X1 U373 ( .A(\u_div/PartRem[18][3] ), .B(\u_div/PartRem[18][2] ), .Y(
        \u_div/SumTmp[17][3] ) );
  OR2X1 U374 ( .A(\u_div/PartRem[17][5] ), .B(\u_div/u_add_PartRem_2_16/n2 ), 
        .Y(\u_div/CryTmp[16][6] ) );
  XNOR2X1 U375 ( .A(\u_div/PartRem[17][3] ), .B(\u_div/PartRem[17][2] ), .Y(
        \u_div/SumTmp[16][3] ) );
  OR2X1 U376 ( .A(\u_div/PartRem[17][2] ), .B(\u_div/PartRem[17][3] ), .Y(
        \u_div/u_add_PartRem_2_16/n3 ) );
  XNOR2X1 U377 ( .A(\u_div/PartRem[16][3] ), .B(\u_div/PartRem[16][2] ), .Y(
        \u_div/SumTmp[15][3] ) );
  OR2X1 U378 ( .A(\u_div/PartRem[15][5] ), .B(\u_div/u_add_PartRem_2_14/n2 ), 
        .Y(\u_div/CryTmp[14][6] ) );
  XNOR2X1 U379 ( .A(\u_div/PartRem[15][3] ), .B(\u_div/PartRem[15][2] ), .Y(
        \u_div/SumTmp[14][3] ) );
  OR2X1 U380 ( .A(\u_div/PartRem[15][2] ), .B(\u_div/PartRem[15][3] ), .Y(
        \u_div/u_add_PartRem_2_14/n3 ) );
  XNOR2X1 U381 ( .A(\u_div/PartRem[14][3] ), .B(\u_div/PartRem[14][2] ), .Y(
        \u_div/SumTmp[13][3] ) );
  OR2X1 U382 ( .A(\u_div/PartRem[13][5] ), .B(\u_div/u_add_PartRem_2_12/n2 ), 
        .Y(\u_div/CryTmp[12][6] ) );
  XNOR2X1 U383 ( .A(\u_div/PartRem[13][3] ), .B(\u_div/PartRem[13][2] ), .Y(
        \u_div/SumTmp[12][3] ) );
  OR2X1 U384 ( .A(\u_div/PartRem[13][2] ), .B(\u_div/PartRem[13][3] ), .Y(
        \u_div/u_add_PartRem_2_12/n3 ) );
  OR2X1 U385 ( .A(\u_div/PartRem[12][5] ), .B(\u_div/u_add_PartRem_2_11/n2 ), 
        .Y(\u_div/CryTmp[11][6] ) );
  XNOR2X1 U386 ( .A(\u_div/PartRem[12][3] ), .B(\u_div/PartRem[12][2] ), .Y(
        \u_div/SumTmp[11][3] ) );
  OR2X1 U387 ( .A(\u_div/PartRem[11][5] ), .B(\u_div/u_add_PartRem_2_10/n2 ), 
        .Y(\u_div/CryTmp[10][6] ) );
  XNOR2X1 U388 ( .A(\u_div/PartRem[11][3] ), .B(\u_div/PartRem[11][2] ), .Y(
        \u_div/SumTmp[10][3] ) );
  OR2X1 U389 ( .A(\u_div/PartRem[10][5] ), .B(\u_div/u_add_PartRem_2_9/n2 ), 
        .Y(\u_div/CryTmp[9][6] ) );
  XNOR2X1 U390 ( .A(\u_div/PartRem[10][3] ), .B(\u_div/PartRem[10][2] ), .Y(
        \u_div/SumTmp[9][3] ) );
  OR2X1 U391 ( .A(\u_div/PartRem[9][5] ), .B(\u_div/u_add_PartRem_2_8/n2 ), 
        .Y(\u_div/CryTmp[8][6] ) );
  XNOR2X1 U392 ( .A(\u_div/PartRem[9][3] ), .B(\u_div/PartRem[9][2] ), .Y(
        \u_div/SumTmp[8][3] ) );
  OR2X1 U393 ( .A(\u_div/PartRem[8][5] ), .B(\u_div/u_add_PartRem_2_7/n2 ), 
        .Y(\u_div/CryTmp[7][6] ) );
  XNOR2X1 U394 ( .A(\u_div/PartRem[8][3] ), .B(\u_div/PartRem[8][2] ), .Y(
        \u_div/SumTmp[7][3] ) );
  OR2X1 U395 ( .A(\u_div/PartRem[7][5] ), .B(\u_div/u_add_PartRem_2_6/n2 ), 
        .Y(\u_div/CryTmp[6][6] ) );
  XNOR2X1 U396 ( .A(\u_div/PartRem[7][3] ), .B(\u_div/PartRem[7][2] ), .Y(
        \u_div/SumTmp[6][3] ) );
  OR2X1 U397 ( .A(\u_div/PartRem[6][5] ), .B(\u_div/u_add_PartRem_2_5/n2 ), 
        .Y(\u_div/CryTmp[5][6] ) );
  XNOR2X1 U398 ( .A(\u_div/PartRem[6][3] ), .B(\u_div/PartRem[6][2] ), .Y(
        \u_div/SumTmp[5][3] ) );
  OR2X1 U399 ( .A(\u_div/PartRem[5][5] ), .B(\u_div/u_add_PartRem_2_4/n2 ), 
        .Y(\u_div/CryTmp[4][6] ) );
  XNOR2X1 U400 ( .A(\u_div/PartRem[5][3] ), .B(\u_div/PartRem[5][2] ), .Y(
        \u_div/SumTmp[4][3] ) );
  OR2X1 U401 ( .A(\u_div/PartRem[4][5] ), .B(\u_div/u_add_PartRem_2_3/n2 ), 
        .Y(\u_div/CryTmp[3][6] ) );
  XNOR2X1 U402 ( .A(\u_div/PartRem[4][3] ), .B(\u_div/PartRem[4][2] ), .Y(
        \u_div/SumTmp[3][3] ) );
  OR2X1 U403 ( .A(\u_div/PartRem[3][5] ), .B(\u_div/u_add_PartRem_2_2/n2 ), 
        .Y(\u_div/CryTmp[2][6] ) );
  XNOR2X1 U404 ( .A(\u_div/PartRem[3][3] ), .B(\u_div/PartRem[3][2] ), .Y(
        \u_div/SumTmp[2][3] ) );
  OR2X1 U405 ( .A(\u_div/PartRem[2][5] ), .B(\u_div/u_add_PartRem_2_1/n2 ), 
        .Y(\u_div/CryTmp[1][6] ) );
  XNOR2X1 U406 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/PartRem[2][2] ), .Y(
        \u_div/SumTmp[1][3] ) );
  NAND2BX1 U407 ( .AN(\u_div/PartRem[1][3] ), .B(n1), .Y(n6) );
  XNOR2X1 U408 ( .A(\u_div/PartRem[63][0] ), .B(\u_div/PartRem[62][0] ), .Y(
        \u_div/SumTmp[59][3] ) );
  XOR2X1 U409 ( .A(\u_div/CryTmp[5][6] ), .B(n4), .Y(\u_div/QInv[5] ) );
  XOR2X1 U410 ( .A(\u_div/CryTmp[57][6] ), .B(n4), .Y(\u_div/QInv[57] ) );
  XOR2X1 U411 ( .A(\u_div/CryTmp[55][6] ), .B(n5), .Y(\u_div/QInv[55] ) );
  XOR2X1 U412 ( .A(\u_div/CryTmp[54][6] ), .B(n4), .Y(\u_div/QInv[54] ) );
  XOR2X1 U413 ( .A(\u_div/CryTmp[44][6] ), .B(n5), .Y(\u_div/QInv[44] ) );
  XOR2X1 U414 ( .A(\u_div/CryTmp[43][6] ), .B(n4), .Y(\u_div/QInv[43] ) );
  XOR2X1 U415 ( .A(\u_div/CryTmp[31][6] ), .B(n5), .Y(\u_div/QInv[31] ) );
  XOR2X1 U416 ( .A(\u_div/CryTmp[18][6] ), .B(n5), .Y(\u_div/QInv[18] ) );
  XOR2X1 U417 ( .A(\u_div/CryTmp[17][6] ), .B(n4), .Y(\u_div/QInv[17] ) );
  XOR2X1 U418 ( .A(\u_div/CryTmp[13][6] ), .B(n4), .Y(\u_div/QInv[13] ) );
  XOR2X1 U419 ( .A(\u_div/CryTmp[0][6] ), .B(n5), .Y(\u_div/QInv[0] ) );
endmodule


module GSIM_DW01_inc_5 ( A, SUM );
  input [63:0] A;
  output [63:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;

  XOR2X1 U2 ( .A(A[63]), .B(n20), .Y(SUM[63]) );
  XNOR2XL U3 ( .A(A[61]), .B(n23), .Y(SUM[61]) );
  NOR3BX1 U4 ( .AN(A[59]), .B(n1), .C(n24), .Y(n22) );
  NOR3BX1 U5 ( .AN(A[55]), .B(n2), .C(n30), .Y(n28) );
  NOR3BX1 U6 ( .AN(A[51]), .B(n3), .C(n34), .Y(n32) );
  NOR3BX1 U7 ( .AN(A[47]), .B(n4), .C(n38), .Y(n36) );
  NOR3BX1 U8 ( .AN(A[43]), .B(n5), .C(n42), .Y(n40) );
  NOR3BX1 U9 ( .AN(A[39]), .B(n6), .C(n46), .Y(n44) );
  NOR3BX1 U10 ( .AN(A[35]), .B(n7), .C(n52), .Y(n50) );
  NOR3BX1 U11 ( .AN(A[31]), .B(n8), .C(n56), .Y(n54) );
  NOR3BX1 U12 ( .AN(A[27]), .B(n9), .C(n60), .Y(n58) );
  NOR3BX1 U13 ( .AN(A[23]), .B(n10), .C(n64), .Y(n62) );
  CLKINVX1 U14 ( .A(A[58]), .Y(n1) );
  CLKINVX1 U15 ( .A(A[54]), .Y(n2) );
  CLKINVX1 U16 ( .A(A[50]), .Y(n3) );
  CLKINVX1 U17 ( .A(A[46]), .Y(n4) );
  CLKINVX1 U18 ( .A(A[42]), .Y(n5) );
  CLKINVX1 U19 ( .A(A[38]), .Y(n6) );
  CLKINVX1 U20 ( .A(A[34]), .Y(n7) );
  CLKINVX1 U21 ( .A(A[30]), .Y(n8) );
  CLKINVX1 U22 ( .A(A[26]), .Y(n9) );
  NOR2BX1 U23 ( .AN(A[62]), .B(n21), .Y(n20) );
  NOR3BX1 U24 ( .AN(A[19]), .B(n11), .C(n68), .Y(n66) );
  NOR3BX1 U25 ( .AN(A[15]), .B(n12), .C(n72), .Y(n70) );
  NOR3BX1 U26 ( .AN(A[11]), .B(n13), .C(n76), .Y(n74) );
  NOR3BX1 U27 ( .AN(A[7]), .B(n14), .C(n19), .Y(n17) );
  NAND3X1 U28 ( .A(A[4]), .B(n26), .C(A[5]), .Y(n19) );
  CLKINVX1 U29 ( .A(A[22]), .Y(n10) );
  CLKINVX1 U30 ( .A(A[18]), .Y(n11) );
  CLKINVX1 U31 ( .A(A[14]), .Y(n12) );
  CLKINVX1 U32 ( .A(A[10]), .Y(n13) );
  CLKINVX1 U33 ( .A(A[6]), .Y(n14) );
  NOR3BX1 U34 ( .AN(A[3]), .B(n15), .C(n48), .Y(n26) );
  NOR2XL U35 ( .A(n24), .B(n1), .Y(n27) );
  NAND2XL U36 ( .A(A[56]), .B(n28), .Y(n29) );
  NOR2XL U37 ( .A(n30), .B(n2), .Y(n31) );
  NAND2XL U38 ( .A(A[52]), .B(n32), .Y(n33) );
  NOR2XL U39 ( .A(n34), .B(n3), .Y(n35) );
  NAND2XL U40 ( .A(A[48]), .B(n36), .Y(n37) );
  NOR2XL U41 ( .A(n38), .B(n4), .Y(n39) );
  NAND2XL U42 ( .A(A[44]), .B(n40), .Y(n41) );
  NOR2XL U43 ( .A(n42), .B(n5), .Y(n43) );
  NAND2XL U44 ( .A(A[40]), .B(n44), .Y(n45) );
  NOR2XL U45 ( .A(n46), .B(n6), .Y(n49) );
  NAND2XL U46 ( .A(A[36]), .B(n50), .Y(n51) );
  NOR2XL U47 ( .A(n52), .B(n7), .Y(n53) );
  NAND2XL U48 ( .A(A[32]), .B(n54), .Y(n55) );
  NOR2XL U49 ( .A(n56), .B(n8), .Y(n57) );
  NAND2XL U50 ( .A(A[28]), .B(n58), .Y(n59) );
  NOR2XL U51 ( .A(n60), .B(n9), .Y(n61) );
  NAND2XL U52 ( .A(A[24]), .B(n62), .Y(n63) );
  NOR2XL U53 ( .A(n64), .B(n10), .Y(n65) );
  NAND2XL U54 ( .A(A[20]), .B(n66), .Y(n67) );
  NOR2XL U55 ( .A(n68), .B(n11), .Y(n69) );
  NAND2XL U56 ( .A(A[16]), .B(n70), .Y(n71) );
  NOR2XL U57 ( .A(n72), .B(n12), .Y(n73) );
  NAND2XL U58 ( .A(A[12]), .B(n74), .Y(n75) );
  NOR2XL U59 ( .A(n76), .B(n13), .Y(n77) );
  NAND2XL U60 ( .A(A[8]), .B(n17), .Y(n16) );
  NOR2XL U61 ( .A(n19), .B(n14), .Y(n18) );
  XOR2XL U62 ( .A(A[60]), .B(n22), .Y(SUM[60]) );
  NAND2XL U63 ( .A(A[60]), .B(n22), .Y(n23) );
  XOR2XL U64 ( .A(n2), .B(n30), .Y(SUM[54]) );
  XNOR2XL U65 ( .A(A[49]), .B(n37), .Y(SUM[49]) );
  XOR2XL U66 ( .A(A[44]), .B(n40), .Y(SUM[44]) );
  XOR2XL U67 ( .A(A[39]), .B(n49), .Y(SUM[39]) );
  XOR2XL U68 ( .A(n7), .B(n52), .Y(SUM[34]) );
  XNOR2XL U69 ( .A(A[29]), .B(n59), .Y(SUM[29]) );
  XOR2XL U70 ( .A(A[24]), .B(n62), .Y(SUM[24]) );
  XNOR2XL U71 ( .A(A[62]), .B(n21), .Y(SUM[62]) );
  NOR2XL U72 ( .A(n48), .B(n15), .Y(n47) );
  CLKINVX1 U73 ( .A(A[2]), .Y(n15) );
  XNOR2X1 U74 ( .A(A[9]), .B(n16), .Y(SUM[9]) );
  XOR2X1 U75 ( .A(A[8]), .B(n17), .Y(SUM[8]) );
  XOR2X1 U76 ( .A(A[7]), .B(n18), .Y(SUM[7]) );
  XOR2X1 U77 ( .A(n14), .B(n19), .Y(SUM[6]) );
  NAND3X1 U78 ( .A(A[60]), .B(n22), .C(A[61]), .Y(n21) );
  XNOR2X1 U79 ( .A(A[5]), .B(n25), .Y(SUM[5]) );
  NAND2X1 U80 ( .A(A[4]), .B(n26), .Y(n25) );
  XOR2X1 U81 ( .A(A[59]), .B(n27), .Y(SUM[59]) );
  XOR2X1 U82 ( .A(n1), .B(n24), .Y(SUM[58]) );
  NAND3X1 U83 ( .A(A[56]), .B(n28), .C(A[57]), .Y(n24) );
  XNOR2X1 U84 ( .A(A[57]), .B(n29), .Y(SUM[57]) );
  XOR2X1 U85 ( .A(A[56]), .B(n28), .Y(SUM[56]) );
  XOR2X1 U86 ( .A(A[55]), .B(n31), .Y(SUM[55]) );
  NAND3X1 U87 ( .A(A[52]), .B(n32), .C(A[53]), .Y(n30) );
  XNOR2X1 U88 ( .A(A[53]), .B(n33), .Y(SUM[53]) );
  XOR2X1 U89 ( .A(A[52]), .B(n32), .Y(SUM[52]) );
  XOR2X1 U90 ( .A(A[51]), .B(n35), .Y(SUM[51]) );
  XOR2X1 U91 ( .A(n3), .B(n34), .Y(SUM[50]) );
  NAND3X1 U92 ( .A(A[48]), .B(n36), .C(A[49]), .Y(n34) );
  XOR2X1 U93 ( .A(A[4]), .B(n26), .Y(SUM[4]) );
  XOR2X1 U94 ( .A(A[48]), .B(n36), .Y(SUM[48]) );
  XOR2X1 U95 ( .A(A[47]), .B(n39), .Y(SUM[47]) );
  XOR2X1 U96 ( .A(n4), .B(n38), .Y(SUM[46]) );
  NAND3X1 U97 ( .A(A[44]), .B(n40), .C(A[45]), .Y(n38) );
  XNOR2X1 U98 ( .A(A[45]), .B(n41), .Y(SUM[45]) );
  XOR2X1 U99 ( .A(A[43]), .B(n43), .Y(SUM[43]) );
  XOR2X1 U100 ( .A(n5), .B(n42), .Y(SUM[42]) );
  NAND3X1 U101 ( .A(A[40]), .B(n44), .C(A[41]), .Y(n42) );
  XNOR2X1 U102 ( .A(A[41]), .B(n45), .Y(SUM[41]) );
  XOR2X1 U103 ( .A(A[40]), .B(n44), .Y(SUM[40]) );
  XOR2X1 U104 ( .A(A[3]), .B(n47), .Y(SUM[3]) );
  XOR2X1 U105 ( .A(n6), .B(n46), .Y(SUM[38]) );
  NAND3X1 U106 ( .A(A[36]), .B(n50), .C(A[37]), .Y(n46) );
  XNOR2X1 U107 ( .A(A[37]), .B(n51), .Y(SUM[37]) );
  XOR2X1 U108 ( .A(A[36]), .B(n50), .Y(SUM[36]) );
  XOR2X1 U109 ( .A(A[35]), .B(n53), .Y(SUM[35]) );
  NAND3X1 U110 ( .A(A[32]), .B(n54), .C(A[33]), .Y(n52) );
  XNOR2X1 U111 ( .A(A[33]), .B(n55), .Y(SUM[33]) );
  XOR2X1 U112 ( .A(A[32]), .B(n54), .Y(SUM[32]) );
  XOR2X1 U113 ( .A(A[31]), .B(n57), .Y(SUM[31]) );
  XOR2X1 U114 ( .A(n8), .B(n56), .Y(SUM[30]) );
  NAND3X1 U115 ( .A(A[28]), .B(n58), .C(A[29]), .Y(n56) );
  XOR2X1 U116 ( .A(n15), .B(n48), .Y(SUM[2]) );
  XOR2X1 U117 ( .A(A[28]), .B(n58), .Y(SUM[28]) );
  XOR2X1 U118 ( .A(A[27]), .B(n61), .Y(SUM[27]) );
  XOR2X1 U119 ( .A(n9), .B(n60), .Y(SUM[26]) );
  NAND3X1 U120 ( .A(A[24]), .B(n62), .C(A[25]), .Y(n60) );
  XNOR2X1 U121 ( .A(A[25]), .B(n63), .Y(SUM[25]) );
  XOR2X1 U122 ( .A(A[23]), .B(n65), .Y(SUM[23]) );
  XOR2X1 U123 ( .A(n10), .B(n64), .Y(SUM[22]) );
  NAND3X1 U124 ( .A(A[20]), .B(n66), .C(A[21]), .Y(n64) );
  XNOR2X1 U125 ( .A(A[21]), .B(n67), .Y(SUM[21]) );
  XOR2X1 U126 ( .A(A[20]), .B(n66), .Y(SUM[20]) );
  XOR2X1 U127 ( .A(A[19]), .B(n69), .Y(SUM[19]) );
  XOR2X1 U128 ( .A(n11), .B(n68), .Y(SUM[18]) );
  NAND3X1 U129 ( .A(A[16]), .B(n70), .C(A[17]), .Y(n68) );
  XNOR2X1 U130 ( .A(A[17]), .B(n71), .Y(SUM[17]) );
  XOR2X1 U131 ( .A(A[16]), .B(n70), .Y(SUM[16]) );
  XOR2X1 U132 ( .A(A[15]), .B(n73), .Y(SUM[15]) );
  XOR2X1 U133 ( .A(n12), .B(n72), .Y(SUM[14]) );
  NAND3X1 U134 ( .A(A[12]), .B(n74), .C(A[13]), .Y(n72) );
  XNOR2X1 U135 ( .A(A[13]), .B(n75), .Y(SUM[13]) );
  XOR2X1 U136 ( .A(A[12]), .B(n74), .Y(SUM[12]) );
  XOR2X1 U137 ( .A(A[11]), .B(n77), .Y(SUM[11]) );
  XOR2X1 U138 ( .A(n13), .B(n76), .Y(SUM[10]) );
  NAND3X1 U139 ( .A(A[8]), .B(n17), .C(A[9]), .Y(n76) );
  NAND2X1 U140 ( .A(A[1]), .B(A[0]), .Y(n48) );
endmodule


module GSIM_DW01_absval_3 ( A, ABSVAL );
  input [63:0] A;
  output [63:0] ABSVAL;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69;
  wire   [63:0] AMUX1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  GSIM_DW01_inc_5 NEG ( .A({n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
        n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
        n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
        n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, 
        n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69}), .SUM({
        AMUX1[63:2], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1}) );
  CLKMX2X2 U1 ( .A(A[61]), .B(AMUX1[61]), .S0(n4), .Y(ABSVAL[61]) );
  CLKINVX1 U2 ( .A(A[60]), .Y(n9) );
  CLKINVX1 U3 ( .A(A[56]), .Y(n13) );
  CLKINVX1 U4 ( .A(A[58]), .Y(n11) );
  CLKINVX1 U5 ( .A(A[54]), .Y(n15) );
  CLKINVX1 U6 ( .A(A[52]), .Y(n17) );
  CLKINVX1 U7 ( .A(A[50]), .Y(n19) );
  CLKINVX1 U8 ( .A(A[48]), .Y(n21) );
  CLKINVX1 U9 ( .A(A[44]), .Y(n25) );
  CLKINVX1 U10 ( .A(A[46]), .Y(n23) );
  CLKINVX1 U11 ( .A(A[42]), .Y(n27) );
  CLKINVX1 U12 ( .A(A[40]), .Y(n29) );
  CLKINVX1 U13 ( .A(A[38]), .Y(n31) );
  CLKINVX1 U14 ( .A(A[36]), .Y(n33) );
  CLKINVX1 U15 ( .A(A[32]), .Y(n37) );
  CLKINVX1 U16 ( .A(A[34]), .Y(n35) );
  CLKINVX1 U17 ( .A(A[30]), .Y(n39) );
  CLKINVX1 U18 ( .A(A[28]), .Y(n41) );
  CLKINVX1 U19 ( .A(A[26]), .Y(n43) );
  CLKINVX1 U20 ( .A(A[24]), .Y(n45) );
  CLKINVX1 U21 ( .A(A[20]), .Y(n49) );
  CLKINVX1 U22 ( .A(A[22]), .Y(n47) );
  CLKINVX1 U23 ( .A(A[18]), .Y(n51) );
  CLKINVX1 U24 ( .A(A[16]), .Y(n53) );
  CLKINVX1 U25 ( .A(A[12]), .Y(n57) );
  CLKINVX1 U26 ( .A(A[14]), .Y(n55) );
  CLKINVX1 U27 ( .A(A[8]), .Y(n61) );
  CLKINVX1 U28 ( .A(A[10]), .Y(n59) );
  CLKINVX1 U29 ( .A(A[6]), .Y(n63) );
  CLKINVX1 U30 ( .A(A[4]), .Y(n65) );
  CLKBUFX2 U31 ( .A(n6), .Y(n5) );
  INVX3 U32 ( .A(n6), .Y(n4) );
  INVX3 U33 ( .A(n5), .Y(n3) );
  INVX3 U34 ( .A(n5), .Y(n2) );
  INVX3 U35 ( .A(n5), .Y(n1) );
  CLKINVX1 U36 ( .A(A[63]), .Y(n6) );
  CLKINVX1 U37 ( .A(A[3]), .Y(n66) );
  CLKINVX1 U38 ( .A(A[2]), .Y(n67) );
  CLKINVX1 U39 ( .A(A[9]), .Y(n60) );
  CLKINVX1 U40 ( .A(A[5]), .Y(n64) );
  CLKINVX1 U41 ( .A(A[19]), .Y(n50) );
  CLKINVX1 U42 ( .A(A[11]), .Y(n58) );
  CLKINVX1 U43 ( .A(A[7]), .Y(n62) );
  CLKINVX1 U44 ( .A(A[21]), .Y(n48) );
  CLKINVX1 U45 ( .A(A[17]), .Y(n52) );
  CLKINVX1 U46 ( .A(A[13]), .Y(n56) );
  CLKINVX1 U47 ( .A(A[51]), .Y(n18) );
  CLKINVX1 U48 ( .A(A[39]), .Y(n30) );
  CLKINVX1 U49 ( .A(A[35]), .Y(n34) );
  CLKINVX1 U50 ( .A(A[31]), .Y(n38) );
  CLKINVX1 U51 ( .A(A[27]), .Y(n42) );
  CLKINVX1 U52 ( .A(A[23]), .Y(n46) );
  CLKINVX1 U53 ( .A(A[15]), .Y(n54) );
  CLKINVX1 U54 ( .A(A[61]), .Y(n8) );
  CLKINVX1 U55 ( .A(A[57]), .Y(n12) );
  CLKINVX1 U56 ( .A(A[53]), .Y(n16) );
  CLKINVX1 U57 ( .A(A[49]), .Y(n20) );
  CLKINVX1 U58 ( .A(A[45]), .Y(n24) );
  CLKINVX1 U59 ( .A(A[41]), .Y(n28) );
  CLKINVX1 U60 ( .A(A[37]), .Y(n32) );
  CLKINVX1 U61 ( .A(A[33]), .Y(n36) );
  CLKINVX1 U62 ( .A(A[29]), .Y(n40) );
  CLKINVX1 U63 ( .A(A[25]), .Y(n44) );
  CLKINVX1 U64 ( .A(A[62]), .Y(n7) );
  CLKINVX1 U65 ( .A(A[59]), .Y(n10) );
  CLKINVX1 U66 ( .A(A[55]), .Y(n14) );
  CLKINVX1 U67 ( .A(A[47]), .Y(n22) );
  CLKINVX1 U68 ( .A(A[43]), .Y(n26) );
  CLKINVX1 U69 ( .A(A[0]), .Y(n69) );
  CLKINVX1 U70 ( .A(A[1]), .Y(n68) );
  CLKMX2X2 U71 ( .A(A[9]), .B(AMUX1[9]), .S0(n3), .Y(ABSVAL[9]) );
  CLKMX2X2 U72 ( .A(A[8]), .B(AMUX1[8]), .S0(n4), .Y(ABSVAL[8]) );
  CLKMX2X2 U73 ( .A(A[7]), .B(AMUX1[7]), .S0(n4), .Y(ABSVAL[7]) );
  CLKMX2X2 U74 ( .A(A[6]), .B(AMUX1[6]), .S0(n4), .Y(ABSVAL[6]) );
  AND2X1 U75 ( .A(AMUX1[63]), .B(n4), .Y(ABSVAL[63]) );
  CLKMX2X2 U76 ( .A(A[62]), .B(AMUX1[62]), .S0(n4), .Y(ABSVAL[62]) );
  CLKMX2X2 U77 ( .A(A[60]), .B(AMUX1[60]), .S0(n4), .Y(ABSVAL[60]) );
  CLKMX2X2 U78 ( .A(A[5]), .B(AMUX1[5]), .S0(n4), .Y(ABSVAL[5]) );
  CLKMX2X2 U79 ( .A(A[59]), .B(AMUX1[59]), .S0(n4), .Y(ABSVAL[59]) );
  CLKMX2X2 U80 ( .A(A[58]), .B(AMUX1[58]), .S0(n4), .Y(ABSVAL[58]) );
  CLKMX2X2 U81 ( .A(A[57]), .B(AMUX1[57]), .S0(n4), .Y(ABSVAL[57]) );
  CLKMX2X2 U82 ( .A(A[56]), .B(AMUX1[56]), .S0(n3), .Y(ABSVAL[56]) );
  CLKMX2X2 U83 ( .A(A[55]), .B(AMUX1[55]), .S0(n3), .Y(ABSVAL[55]) );
  CLKMX2X2 U84 ( .A(A[54]), .B(AMUX1[54]), .S0(n3), .Y(ABSVAL[54]) );
  CLKMX2X2 U85 ( .A(A[53]), .B(AMUX1[53]), .S0(n3), .Y(ABSVAL[53]) );
  CLKMX2X2 U86 ( .A(A[52]), .B(AMUX1[52]), .S0(n3), .Y(ABSVAL[52]) );
  CLKMX2X2 U87 ( .A(A[51]), .B(AMUX1[51]), .S0(n3), .Y(ABSVAL[51]) );
  CLKMX2X2 U88 ( .A(A[50]), .B(AMUX1[50]), .S0(n3), .Y(ABSVAL[50]) );
  CLKMX2X2 U89 ( .A(A[4]), .B(AMUX1[4]), .S0(n3), .Y(ABSVAL[4]) );
  CLKMX2X2 U90 ( .A(A[49]), .B(AMUX1[49]), .S0(n3), .Y(ABSVAL[49]) );
  CLKMX2X2 U91 ( .A(A[48]), .B(AMUX1[48]), .S0(n3), .Y(ABSVAL[48]) );
  CLKMX2X2 U92 ( .A(A[47]), .B(AMUX1[47]), .S0(n3), .Y(ABSVAL[47]) );
  CLKMX2X2 U93 ( .A(A[46]), .B(AMUX1[46]), .S0(n3), .Y(ABSVAL[46]) );
  CLKMX2X2 U94 ( .A(A[45]), .B(AMUX1[45]), .S0(n3), .Y(ABSVAL[45]) );
  CLKMX2X2 U95 ( .A(A[44]), .B(AMUX1[44]), .S0(n2), .Y(ABSVAL[44]) );
  CLKMX2X2 U96 ( .A(A[43]), .B(AMUX1[43]), .S0(n2), .Y(ABSVAL[43]) );
  CLKMX2X2 U97 ( .A(A[42]), .B(AMUX1[42]), .S0(n2), .Y(ABSVAL[42]) );
  CLKMX2X2 U98 ( .A(A[41]), .B(AMUX1[41]), .S0(n2), .Y(ABSVAL[41]) );
  CLKMX2X2 U99 ( .A(A[40]), .B(AMUX1[40]), .S0(n2), .Y(ABSVAL[40]) );
  CLKMX2X2 U100 ( .A(A[3]), .B(AMUX1[3]), .S0(n2), .Y(ABSVAL[3]) );
  CLKMX2X2 U101 ( .A(A[39]), .B(AMUX1[39]), .S0(n2), .Y(ABSVAL[39]) );
  CLKMX2X2 U102 ( .A(A[38]), .B(AMUX1[38]), .S0(n2), .Y(ABSVAL[38]) );
  CLKMX2X2 U103 ( .A(A[37]), .B(AMUX1[37]), .S0(n2), .Y(ABSVAL[37]) );
  CLKMX2X2 U104 ( .A(A[36]), .B(AMUX1[36]), .S0(n2), .Y(ABSVAL[36]) );
  CLKMX2X2 U105 ( .A(A[35]), .B(AMUX1[35]), .S0(n2), .Y(ABSVAL[35]) );
  CLKMX2X2 U106 ( .A(A[34]), .B(AMUX1[34]), .S0(n2), .Y(ABSVAL[34]) );
  CLKMX2X2 U107 ( .A(A[33]), .B(AMUX1[33]), .S0(n1), .Y(ABSVAL[33]) );
  CLKMX2X2 U108 ( .A(A[32]), .B(AMUX1[32]), .S0(n1), .Y(ABSVAL[32]) );
  CLKMX2X2 U109 ( .A(A[31]), .B(AMUX1[31]), .S0(n1), .Y(ABSVAL[31]) );
  CLKMX2X2 U110 ( .A(A[30]), .B(AMUX1[30]), .S0(n1), .Y(ABSVAL[30]) );
  CLKMX2X2 U111 ( .A(A[2]), .B(AMUX1[2]), .S0(n1), .Y(ABSVAL[2]) );
  CLKMX2X2 U112 ( .A(A[29]), .B(AMUX1[29]), .S0(n1), .Y(ABSVAL[29]) );
  CLKMX2X2 U113 ( .A(A[28]), .B(AMUX1[28]), .S0(n1), .Y(ABSVAL[28]) );
  CLKMX2X2 U114 ( .A(A[27]), .B(AMUX1[27]), .S0(n1), .Y(ABSVAL[27]) );
  CLKMX2X2 U115 ( .A(A[26]), .B(AMUX1[26]), .S0(n1), .Y(ABSVAL[26]) );
  CLKMX2X2 U116 ( .A(A[25]), .B(AMUX1[25]), .S0(n1), .Y(ABSVAL[25]) );
  CLKMX2X2 U117 ( .A(A[24]), .B(AMUX1[24]), .S0(n1), .Y(ABSVAL[24]) );
  CLKMX2X2 U118 ( .A(A[23]), .B(AMUX1[23]), .S0(n1), .Y(ABSVAL[23]) );
  CLKMX2X2 U119 ( .A(A[22]), .B(AMUX1[22]), .S0(n1), .Y(ABSVAL[22]) );
  CLKMX2X2 U120 ( .A(A[21]), .B(AMUX1[21]), .S0(n1), .Y(ABSVAL[21]) );
  CLKMX2X2 U121 ( .A(A[20]), .B(AMUX1[20]), .S0(n1), .Y(ABSVAL[20]) );
  CLKMX2X2 U122 ( .A(A[19]), .B(AMUX1[19]), .S0(n1), .Y(ABSVAL[19]) );
  CLKMX2X2 U123 ( .A(A[18]), .B(AMUX1[18]), .S0(n1), .Y(ABSVAL[18]) );
  CLKMX2X2 U124 ( .A(A[17]), .B(AMUX1[17]), .S0(n2), .Y(ABSVAL[17]) );
  CLKMX2X2 U125 ( .A(A[16]), .B(AMUX1[16]), .S0(n2), .Y(ABSVAL[16]) );
  CLKMX2X2 U126 ( .A(A[15]), .B(AMUX1[15]), .S0(n2), .Y(ABSVAL[15]) );
  CLKMX2X2 U127 ( .A(A[14]), .B(AMUX1[14]), .S0(n2), .Y(ABSVAL[14]) );
  CLKMX2X2 U128 ( .A(A[13]), .B(AMUX1[13]), .S0(n3), .Y(ABSVAL[13]) );
  CLKMX2X2 U129 ( .A(A[12]), .B(AMUX1[12]), .S0(n3), .Y(ABSVAL[12]) );
  CLKMX2X2 U130 ( .A(A[11]), .B(AMUX1[11]), .S0(n3), .Y(ABSVAL[11]) );
  CLKMX2X2 U131 ( .A(A[10]), .B(AMUX1[10]), .S0(n2), .Y(ABSVAL[10]) );
endmodule


module GSIM_DW_inc_3 ( carry_in, a, carry_out, sum );
  input [63:0] a;
  output [63:0] sum;
  input carry_in;
  output carry_out;
  wire   \sum[63] , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63;
  assign sum[62] = \sum[63] ;
  assign sum[61] = \sum[63] ;
  assign sum[63] = \sum[63] ;

  ADDHXL U23 ( .A(a[43]), .B(n21), .CO(n20), .S(sum[43]) );
  ADDHXL U25 ( .A(a[41]), .B(n23), .CO(n22), .S(sum[41]) );
  ADDHXL U35 ( .A(a[31]), .B(n33), .CO(n32), .S(sum[31]) );
  ADDHXL U46 ( .A(a[20]), .B(n44), .CO(n43), .S(sum[20]) );
  ADDHXL U50 ( .A(a[16]), .B(n48), .CO(n47), .S(sum[16]) );
  ADDHXL U54 ( .A(a[12]), .B(n52), .CO(n51), .S(sum[12]) );
  ADDHXL U56 ( .A(a[10]), .B(n54), .CO(n53), .S(sum[10]) );
  ADDHXL U60 ( .A(a[6]), .B(n58), .CO(n57), .S(sum[6]) );
  ADDHXL U62 ( .A(a[4]), .B(n60), .CO(n59), .S(sum[4]) );
  ADDHXL U66 ( .A(carry_in), .B(a[0]), .CO(n63), .S(sum[0]) );
  ADDHXL U70 ( .A(a[13]), .B(n51), .CO(n50), .S(sum[13]) );
  ADDHXL U71 ( .A(a[17]), .B(n47), .CO(n46), .S(sum[17]) );
  ADDHXL U72 ( .A(a[23]), .B(n41), .CO(n40), .S(sum[23]) );
  ADDHXL U73 ( .A(a[21]), .B(n43), .CO(n42), .S(sum[21]) );
  ADDHXL U74 ( .A(a[9]), .B(n55), .CO(n54), .S(sum[9]) );
  ADDHXL U75 ( .A(a[3]), .B(n61), .CO(n60), .S(sum[3]) );
  ADDHXL U76 ( .A(a[7]), .B(n57), .CO(n56), .S(sum[7]) );
  ADDHXL U77 ( .A(a[26]), .B(n38), .CO(n37), .S(sum[26]) );
  ADDHXL U78 ( .A(a[29]), .B(n35), .CO(n34), .S(sum[29]) );
  ADDHXL U79 ( .A(a[32]), .B(n32), .CO(n31), .S(sum[32]) );
  ADDHXL U80 ( .A(a[35]), .B(n29), .CO(n28), .S(sum[35]) );
  ADDHXL U81 ( .A(a[39]), .B(n25), .CO(n24), .S(sum[39]) );
  ADDHXL U82 ( .A(a[42]), .B(n22), .CO(n21), .S(sum[42]) );
  ADDHXL U83 ( .A(a[46]), .B(n18), .CO(n17), .S(sum[46]) );
  ADDHXL U84 ( .A(a[50]), .B(n14), .CO(n13), .S(sum[50]) );
  ADDHXL U85 ( .A(a[55]), .B(n9), .CO(n8), .S(sum[55]) );
  ADDHXL U86 ( .A(a[58]), .B(n6), .CO(n5), .S(sum[58]) );
  ADDHXL U87 ( .A(a[45]), .B(n19), .CO(n18), .S(sum[45]) );
  ADDHXL U88 ( .A(a[44]), .B(n20), .CO(n19), .S(sum[44]) );
  ADDHX1 U89 ( .A(a[11]), .B(n53), .CO(n52), .S(sum[11]) );
  ADDHX1 U90 ( .A(a[5]), .B(n59), .CO(n58), .S(sum[5]) );
  ADDHX1 U91 ( .A(a[48]), .B(n16), .CO(n15), .S(sum[48]) );
  ADDHX1 U92 ( .A(a[56]), .B(n8), .CO(n7), .S(sum[56]) );
  ADDHX1 U93 ( .A(a[37]), .B(n27), .CO(n26), .S(sum[37]) );
  ADDHX1 U94 ( .A(a[53]), .B(n11), .CO(n10), .S(sum[53]) );
  ADDHX1 U95 ( .A(a[19]), .B(n45), .CO(n44), .S(sum[19]) );
  ADDHX1 U96 ( .A(a[1]), .B(n63), .CO(n62), .S(sum[1]) );
  ADDHX1 U97 ( .A(a[34]), .B(n30), .CO(n29), .S(sum[34]) );
  ADDHX1 U98 ( .A(a[15]), .B(n49), .CO(n48), .S(sum[15]) );
  ADDHXL U99 ( .A(a[51]), .B(n13), .CO(n12), .S(sum[51]) );
  ADDHXL U100 ( .A(a[30]), .B(n34), .CO(n33), .S(sum[30]) );
  ADDHXL U101 ( .A(a[40]), .B(n24), .CO(n23), .S(sum[40]) );
  ADDHXL U102 ( .A(a[24]), .B(n40), .CO(n39), .S(sum[24]) );
  ADDHXL U103 ( .A(a[27]), .B(n37), .CO(n36), .S(sum[27]) );
  NOR2BX1 U104 ( .AN(a[60]), .B(n4), .Y(\sum[63] ) );
  XOR2XL U105 ( .A(n4), .B(a[60]), .Y(sum[60]) );
  ADDHXL U106 ( .A(a[54]), .B(n10), .CO(n9), .S(sum[54]) );
  ADDHXL U107 ( .A(a[25]), .B(n39), .CO(n38), .S(sum[25]) );
  ADDHXL U108 ( .A(a[57]), .B(n7), .CO(n6), .S(sum[57]) );
  ADDHXL U109 ( .A(a[59]), .B(n5), .CO(n4), .S(sum[59]) );
  ADDHXL U110 ( .A(a[52]), .B(n12), .CO(n11), .S(sum[52]) );
  ADDHXL U111 ( .A(a[14]), .B(n50), .CO(n49), .S(sum[14]) );
  ADDHXL U112 ( .A(a[22]), .B(n42), .CO(n41), .S(sum[22]) );
  ADDHXL U113 ( .A(a[33]), .B(n31), .CO(n30), .S(sum[33]) );
  ADDHXL U114 ( .A(a[2]), .B(n62), .CO(n61), .S(sum[2]) );
  ADDHXL U115 ( .A(a[49]), .B(n15), .CO(n14), .S(sum[49]) );
  ADDHXL U116 ( .A(a[36]), .B(n28), .CO(n27), .S(sum[36]) );
  ADDHXL U117 ( .A(a[47]), .B(n17), .CO(n16), .S(sum[47]) );
  ADDHXL U118 ( .A(a[8]), .B(n56), .CO(n55), .S(sum[8]) );
  ADDHXL U119 ( .A(a[18]), .B(n46), .CO(n45), .S(sum[18]) );
  ADDHXL U120 ( .A(a[28]), .B(n36), .CO(n35), .S(sum[28]) );
  ADDHXL U121 ( .A(a[38]), .B(n26), .CO(n25), .S(sum[38]) );
endmodule


module GSIM_DW_div_tc_3 ( a, b, quotient, remainder, divide_by_0 );
  input [63:0] a;
  input [5:0] b;
  output [63:0] quotient;
  output [5:0] remainder;
  output divide_by_0;
  wire   \u_div/QInv[63] , \u_div/QInv[59] , \u_div/QInv[58] ,
         \u_div/QInv[57] , \u_div/QInv[56] , \u_div/QInv[55] ,
         \u_div/QInv[54] , \u_div/QInv[53] , \u_div/QInv[52] ,
         \u_div/QInv[51] , \u_div/QInv[50] , \u_div/QInv[49] ,
         \u_div/QInv[48] , \u_div/QInv[47] , \u_div/QInv[46] ,
         \u_div/QInv[45] , \u_div/QInv[44] , \u_div/QInv[43] ,
         \u_div/QInv[42] , \u_div/QInv[41] , \u_div/QInv[40] ,
         \u_div/QInv[39] , \u_div/QInv[38] , \u_div/QInv[37] ,
         \u_div/QInv[36] , \u_div/QInv[35] , \u_div/QInv[34] ,
         \u_div/QInv[33] , \u_div/QInv[32] , \u_div/QInv[31] ,
         \u_div/QInv[30] , \u_div/QInv[29] , \u_div/QInv[28] ,
         \u_div/QInv[27] , \u_div/QInv[26] , \u_div/QInv[25] ,
         \u_div/QInv[24] , \u_div/QInv[23] , \u_div/QInv[22] ,
         \u_div/QInv[21] , \u_div/QInv[20] , \u_div/QInv[19] ,
         \u_div/QInv[18] , \u_div/QInv[17] , \u_div/QInv[16] ,
         \u_div/QInv[15] , \u_div/QInv[14] , \u_div/QInv[13] ,
         \u_div/QInv[12] , \u_div/QInv[11] , \u_div/QInv[10] , \u_div/QInv[9] ,
         \u_div/QInv[8] , \u_div/QInv[7] , \u_div/QInv[6] , \u_div/QInv[5] ,
         \u_div/QInv[4] , \u_div/QInv[3] , \u_div/QInv[2] , \u_div/QInv[1] ,
         \u_div/QInv[0] , \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] ,
         \u_div/SumTmp[1][3] , \u_div/SumTmp[1][4] , \u_div/SumTmp[2][1] ,
         \u_div/SumTmp[2][2] , \u_div/SumTmp[2][3] , \u_div/SumTmp[2][4] ,
         \u_div/SumTmp[3][1] , \u_div/SumTmp[3][2] , \u_div/SumTmp[3][3] ,
         \u_div/SumTmp[3][4] , \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] ,
         \u_div/SumTmp[4][3] , \u_div/SumTmp[4][4] , \u_div/SumTmp[5][1] ,
         \u_div/SumTmp[5][2] , \u_div/SumTmp[5][3] , \u_div/SumTmp[5][4] ,
         \u_div/SumTmp[6][1] , \u_div/SumTmp[6][2] , \u_div/SumTmp[6][3] ,
         \u_div/SumTmp[6][4] , \u_div/SumTmp[7][1] , \u_div/SumTmp[7][2] ,
         \u_div/SumTmp[7][3] , \u_div/SumTmp[7][4] , \u_div/SumTmp[8][1] ,
         \u_div/SumTmp[8][2] , \u_div/SumTmp[8][3] , \u_div/SumTmp[8][4] ,
         \u_div/SumTmp[9][1] , \u_div/SumTmp[9][2] , \u_div/SumTmp[9][3] ,
         \u_div/SumTmp[9][4] , \u_div/SumTmp[10][1] , \u_div/SumTmp[10][2] ,
         \u_div/SumTmp[10][3] , \u_div/SumTmp[10][4] , \u_div/SumTmp[11][1] ,
         \u_div/SumTmp[11][2] , \u_div/SumTmp[11][3] , \u_div/SumTmp[11][4] ,
         \u_div/SumTmp[12][1] , \u_div/SumTmp[12][2] , \u_div/SumTmp[12][3] ,
         \u_div/SumTmp[12][4] , \u_div/SumTmp[13][1] , \u_div/SumTmp[13][2] ,
         \u_div/SumTmp[13][3] , \u_div/SumTmp[13][4] , \u_div/SumTmp[14][1] ,
         \u_div/SumTmp[14][2] , \u_div/SumTmp[14][3] , \u_div/SumTmp[14][4] ,
         \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] , \u_div/SumTmp[15][3] ,
         \u_div/SumTmp[15][4] , \u_div/SumTmp[16][1] , \u_div/SumTmp[16][2] ,
         \u_div/SumTmp[16][3] , \u_div/SumTmp[16][4] , \u_div/SumTmp[17][1] ,
         \u_div/SumTmp[17][2] , \u_div/SumTmp[17][3] , \u_div/SumTmp[17][4] ,
         \u_div/SumTmp[18][1] , \u_div/SumTmp[18][2] , \u_div/SumTmp[18][3] ,
         \u_div/SumTmp[18][4] , \u_div/SumTmp[19][1] , \u_div/SumTmp[19][2] ,
         \u_div/SumTmp[19][3] , \u_div/SumTmp[19][4] , \u_div/SumTmp[20][1] ,
         \u_div/SumTmp[20][2] , \u_div/SumTmp[20][3] , \u_div/SumTmp[20][4] ,
         \u_div/SumTmp[21][1] , \u_div/SumTmp[21][2] , \u_div/SumTmp[21][3] ,
         \u_div/SumTmp[21][4] , \u_div/SumTmp[22][1] , \u_div/SumTmp[22][2] ,
         \u_div/SumTmp[22][3] , \u_div/SumTmp[22][4] , \u_div/SumTmp[23][1] ,
         \u_div/SumTmp[23][2] , \u_div/SumTmp[23][3] , \u_div/SumTmp[23][4] ,
         \u_div/SumTmp[24][1] , \u_div/SumTmp[24][2] , \u_div/SumTmp[24][3] ,
         \u_div/SumTmp[24][4] , \u_div/SumTmp[25][1] , \u_div/SumTmp[25][2] ,
         \u_div/SumTmp[25][3] , \u_div/SumTmp[25][4] , \u_div/SumTmp[26][1] ,
         \u_div/SumTmp[26][2] , \u_div/SumTmp[26][3] , \u_div/SumTmp[26][4] ,
         \u_div/SumTmp[27][1] , \u_div/SumTmp[27][2] , \u_div/SumTmp[27][3] ,
         \u_div/SumTmp[27][4] , \u_div/SumTmp[28][1] , \u_div/SumTmp[28][2] ,
         \u_div/SumTmp[28][3] , \u_div/SumTmp[28][4] , \u_div/SumTmp[29][1] ,
         \u_div/SumTmp[29][2] , \u_div/SumTmp[29][3] , \u_div/SumTmp[29][4] ,
         \u_div/SumTmp[30][1] , \u_div/SumTmp[30][2] , \u_div/SumTmp[30][3] ,
         \u_div/SumTmp[30][4] , \u_div/SumTmp[31][1] , \u_div/SumTmp[31][2] ,
         \u_div/SumTmp[31][3] , \u_div/SumTmp[31][4] , \u_div/SumTmp[32][1] ,
         \u_div/SumTmp[32][2] , \u_div/SumTmp[32][3] , \u_div/SumTmp[32][4] ,
         \u_div/SumTmp[33][1] , \u_div/SumTmp[33][2] , \u_div/SumTmp[33][3] ,
         \u_div/SumTmp[33][4] , \u_div/SumTmp[34][1] , \u_div/SumTmp[34][2] ,
         \u_div/SumTmp[34][3] , \u_div/SumTmp[34][4] , \u_div/SumTmp[35][1] ,
         \u_div/SumTmp[35][2] , \u_div/SumTmp[35][3] , \u_div/SumTmp[35][4] ,
         \u_div/SumTmp[36][1] , \u_div/SumTmp[36][2] , \u_div/SumTmp[36][3] ,
         \u_div/SumTmp[36][4] , \u_div/SumTmp[37][1] , \u_div/SumTmp[37][2] ,
         \u_div/SumTmp[37][3] , \u_div/SumTmp[37][4] , \u_div/SumTmp[38][1] ,
         \u_div/SumTmp[38][2] , \u_div/SumTmp[38][3] , \u_div/SumTmp[38][4] ,
         \u_div/SumTmp[39][1] , \u_div/SumTmp[39][2] , \u_div/SumTmp[39][3] ,
         \u_div/SumTmp[39][4] , \u_div/SumTmp[40][1] , \u_div/SumTmp[40][2] ,
         \u_div/SumTmp[40][3] , \u_div/SumTmp[40][4] , \u_div/SumTmp[41][1] ,
         \u_div/SumTmp[41][2] , \u_div/SumTmp[41][3] , \u_div/SumTmp[41][4] ,
         \u_div/SumTmp[42][1] , \u_div/SumTmp[42][2] , \u_div/SumTmp[42][3] ,
         \u_div/SumTmp[42][4] , \u_div/SumTmp[43][1] , \u_div/SumTmp[43][2] ,
         \u_div/SumTmp[43][3] , \u_div/SumTmp[43][4] , \u_div/SumTmp[44][1] ,
         \u_div/SumTmp[44][2] , \u_div/SumTmp[44][3] , \u_div/SumTmp[44][4] ,
         \u_div/SumTmp[45][1] , \u_div/SumTmp[45][2] , \u_div/SumTmp[45][3] ,
         \u_div/SumTmp[45][4] , \u_div/SumTmp[46][1] , \u_div/SumTmp[46][2] ,
         \u_div/SumTmp[46][3] , \u_div/SumTmp[46][4] , \u_div/SumTmp[47][1] ,
         \u_div/SumTmp[47][2] , \u_div/SumTmp[47][3] , \u_div/SumTmp[47][4] ,
         \u_div/SumTmp[48][1] , \u_div/SumTmp[48][2] , \u_div/SumTmp[48][3] ,
         \u_div/SumTmp[48][4] , \u_div/SumTmp[49][1] , \u_div/SumTmp[49][2] ,
         \u_div/SumTmp[49][3] , \u_div/SumTmp[49][4] , \u_div/SumTmp[50][1] ,
         \u_div/SumTmp[50][2] , \u_div/SumTmp[50][3] , \u_div/SumTmp[50][4] ,
         \u_div/SumTmp[51][1] , \u_div/SumTmp[51][2] , \u_div/SumTmp[51][3] ,
         \u_div/SumTmp[51][4] , \u_div/SumTmp[52][1] , \u_div/SumTmp[52][2] ,
         \u_div/SumTmp[52][3] , \u_div/SumTmp[52][4] , \u_div/SumTmp[53][1] ,
         \u_div/SumTmp[53][2] , \u_div/SumTmp[53][3] , \u_div/SumTmp[53][4] ,
         \u_div/SumTmp[54][1] , \u_div/SumTmp[54][2] , \u_div/SumTmp[54][3] ,
         \u_div/SumTmp[54][4] , \u_div/SumTmp[55][1] , \u_div/SumTmp[55][2] ,
         \u_div/SumTmp[55][3] , \u_div/SumTmp[55][4] , \u_div/SumTmp[56][1] ,
         \u_div/SumTmp[56][2] , \u_div/SumTmp[56][3] , \u_div/SumTmp[56][4] ,
         \u_div/SumTmp[57][1] , \u_div/SumTmp[57][2] , \u_div/SumTmp[57][3] ,
         \u_div/SumTmp[57][4] , \u_div/SumTmp[58][1] , \u_div/SumTmp[58][2] ,
         \u_div/SumTmp[58][3] , \u_div/SumTmp[58][4] , \u_div/SumTmp[59][3] ,
         \u_div/SumTmp[59][4] , \u_div/CryTmp[0][6] , \u_div/CryTmp[1][6] ,
         \u_div/CryTmp[2][6] , \u_div/CryTmp[3][6] , \u_div/CryTmp[4][6] ,
         \u_div/CryTmp[5][6] , \u_div/CryTmp[6][6] , \u_div/CryTmp[7][6] ,
         \u_div/CryTmp[8][6] , \u_div/CryTmp[9][6] , \u_div/CryTmp[10][6] ,
         \u_div/CryTmp[11][6] , \u_div/CryTmp[12][6] , \u_div/CryTmp[13][6] ,
         \u_div/CryTmp[14][6] , \u_div/CryTmp[15][6] , \u_div/CryTmp[16][6] ,
         \u_div/CryTmp[17][6] , \u_div/CryTmp[18][6] , \u_div/CryTmp[19][6] ,
         \u_div/CryTmp[20][6] , \u_div/CryTmp[21][6] , \u_div/CryTmp[22][6] ,
         \u_div/CryTmp[23][6] , \u_div/CryTmp[24][6] , \u_div/CryTmp[25][6] ,
         \u_div/CryTmp[26][6] , \u_div/CryTmp[27][6] , \u_div/CryTmp[28][6] ,
         \u_div/CryTmp[29][6] , \u_div/CryTmp[30][6] , \u_div/CryTmp[31][6] ,
         \u_div/CryTmp[32][6] , \u_div/CryTmp[33][6] , \u_div/CryTmp[34][6] ,
         \u_div/CryTmp[35][6] , \u_div/CryTmp[36][6] , \u_div/CryTmp[37][6] ,
         \u_div/CryTmp[38][6] , \u_div/CryTmp[39][6] , \u_div/CryTmp[40][6] ,
         \u_div/CryTmp[41][6] , \u_div/CryTmp[42][6] , \u_div/CryTmp[43][6] ,
         \u_div/CryTmp[44][6] , \u_div/CryTmp[45][6] , \u_div/CryTmp[46][6] ,
         \u_div/CryTmp[47][6] , \u_div/CryTmp[48][6] , \u_div/CryTmp[49][6] ,
         \u_div/CryTmp[50][6] , \u_div/CryTmp[51][6] , \u_div/CryTmp[52][6] ,
         \u_div/CryTmp[53][6] , \u_div/CryTmp[54][6] , \u_div/CryTmp[55][6] ,
         \u_div/CryTmp[56][6] , \u_div/CryTmp[57][6] , \u_div/CryTmp[58][6] ,
         \u_div/CryTmp[59][6] , \u_div/PartRem[1][3] , \u_div/PartRem[1][4] ,
         \u_div/PartRem[1][5] , \u_div/PartRem[2][2] , \u_div/PartRem[2][3] ,
         \u_div/PartRem[2][4] , \u_div/PartRem[2][5] , \u_div/PartRem[3][0] ,
         \u_div/PartRem[3][2] , \u_div/PartRem[3][3] , \u_div/PartRem[3][4] ,
         \u_div/PartRem[3][5] , \u_div/PartRem[4][0] , \u_div/PartRem[4][2] ,
         \u_div/PartRem[4][3] , \u_div/PartRem[4][4] , \u_div/PartRem[4][5] ,
         \u_div/PartRem[5][0] , \u_div/PartRem[5][2] , \u_div/PartRem[5][3] ,
         \u_div/PartRem[5][4] , \u_div/PartRem[5][5] , \u_div/PartRem[6][0] ,
         \u_div/PartRem[6][2] , \u_div/PartRem[6][3] , \u_div/PartRem[6][4] ,
         \u_div/PartRem[6][5] , \u_div/PartRem[7][0] , \u_div/PartRem[7][2] ,
         \u_div/PartRem[7][3] , \u_div/PartRem[7][4] , \u_div/PartRem[7][5] ,
         \u_div/PartRem[8][0] , \u_div/PartRem[8][2] , \u_div/PartRem[8][3] ,
         \u_div/PartRem[8][4] , \u_div/PartRem[8][5] , \u_div/PartRem[9][0] ,
         \u_div/PartRem[9][2] , \u_div/PartRem[9][3] , \u_div/PartRem[9][4] ,
         \u_div/PartRem[9][5] , \u_div/PartRem[10][0] , \u_div/PartRem[10][2] ,
         \u_div/PartRem[10][3] , \u_div/PartRem[10][4] ,
         \u_div/PartRem[10][5] , \u_div/PartRem[11][0] ,
         \u_div/PartRem[11][2] , \u_div/PartRem[11][3] ,
         \u_div/PartRem[11][4] , \u_div/PartRem[11][5] ,
         \u_div/PartRem[12][0] , \u_div/PartRem[12][2] ,
         \u_div/PartRem[12][3] , \u_div/PartRem[12][4] ,
         \u_div/PartRem[12][5] , \u_div/PartRem[13][0] ,
         \u_div/PartRem[13][2] , \u_div/PartRem[13][3] ,
         \u_div/PartRem[13][4] , \u_div/PartRem[13][5] ,
         \u_div/PartRem[14][0] , \u_div/PartRem[14][2] ,
         \u_div/PartRem[14][3] , \u_div/PartRem[14][4] ,
         \u_div/PartRem[14][5] , \u_div/PartRem[15][0] ,
         \u_div/PartRem[15][2] , \u_div/PartRem[15][3] ,
         \u_div/PartRem[15][4] , \u_div/PartRem[15][5] ,
         \u_div/PartRem[16][0] , \u_div/PartRem[16][2] ,
         \u_div/PartRem[16][3] , \u_div/PartRem[16][4] ,
         \u_div/PartRem[16][5] , \u_div/PartRem[17][0] ,
         \u_div/PartRem[17][2] , \u_div/PartRem[17][3] ,
         \u_div/PartRem[17][4] , \u_div/PartRem[17][5] ,
         \u_div/PartRem[18][0] , \u_div/PartRem[18][2] ,
         \u_div/PartRem[18][3] , \u_div/PartRem[18][4] ,
         \u_div/PartRem[18][5] , \u_div/PartRem[19][0] ,
         \u_div/PartRem[19][2] , \u_div/PartRem[19][3] ,
         \u_div/PartRem[19][4] , \u_div/PartRem[19][5] ,
         \u_div/PartRem[20][0] , \u_div/PartRem[20][2] ,
         \u_div/PartRem[20][3] , \u_div/PartRem[20][4] ,
         \u_div/PartRem[20][5] , \u_div/PartRem[21][0] ,
         \u_div/PartRem[21][2] , \u_div/PartRem[21][3] ,
         \u_div/PartRem[21][4] , \u_div/PartRem[21][5] ,
         \u_div/PartRem[22][0] , \u_div/PartRem[22][2] ,
         \u_div/PartRem[22][3] , \u_div/PartRem[22][4] ,
         \u_div/PartRem[22][5] , \u_div/PartRem[23][0] ,
         \u_div/PartRem[23][2] , \u_div/PartRem[23][3] ,
         \u_div/PartRem[23][4] , \u_div/PartRem[23][5] ,
         \u_div/PartRem[24][0] , \u_div/PartRem[24][2] ,
         \u_div/PartRem[24][3] , \u_div/PartRem[24][4] ,
         \u_div/PartRem[24][5] , \u_div/PartRem[25][0] ,
         \u_div/PartRem[25][2] , \u_div/PartRem[25][3] ,
         \u_div/PartRem[25][4] , \u_div/PartRem[25][5] ,
         \u_div/PartRem[26][0] , \u_div/PartRem[26][2] ,
         \u_div/PartRem[26][3] , \u_div/PartRem[26][4] ,
         \u_div/PartRem[26][5] , \u_div/PartRem[27][0] ,
         \u_div/PartRem[27][2] , \u_div/PartRem[27][3] ,
         \u_div/PartRem[27][4] , \u_div/PartRem[27][5] ,
         \u_div/PartRem[28][0] , \u_div/PartRem[28][2] ,
         \u_div/PartRem[28][3] , \u_div/PartRem[28][4] ,
         \u_div/PartRem[28][5] , \u_div/PartRem[29][0] ,
         \u_div/PartRem[29][2] , \u_div/PartRem[29][3] ,
         \u_div/PartRem[29][4] , \u_div/PartRem[29][5] ,
         \u_div/PartRem[30][0] , \u_div/PartRem[30][2] ,
         \u_div/PartRem[30][3] , \u_div/PartRem[30][4] ,
         \u_div/PartRem[30][5] , \u_div/PartRem[31][0] ,
         \u_div/PartRem[31][2] , \u_div/PartRem[31][3] ,
         \u_div/PartRem[31][4] , \u_div/PartRem[31][5] ,
         \u_div/PartRem[32][0] , \u_div/PartRem[32][2] ,
         \u_div/PartRem[32][3] , \u_div/PartRem[32][4] ,
         \u_div/PartRem[32][5] , \u_div/PartRem[33][0] ,
         \u_div/PartRem[33][2] , \u_div/PartRem[33][3] ,
         \u_div/PartRem[33][4] , \u_div/PartRem[33][5] ,
         \u_div/PartRem[34][0] , \u_div/PartRem[34][2] ,
         \u_div/PartRem[34][3] , \u_div/PartRem[34][4] ,
         \u_div/PartRem[34][5] , \u_div/PartRem[35][0] ,
         \u_div/PartRem[35][2] , \u_div/PartRem[35][3] ,
         \u_div/PartRem[35][4] , \u_div/PartRem[35][5] ,
         \u_div/PartRem[36][0] , \u_div/PartRem[36][2] ,
         \u_div/PartRem[36][3] , \u_div/PartRem[36][4] ,
         \u_div/PartRem[36][5] , \u_div/PartRem[37][0] ,
         \u_div/PartRem[37][2] , \u_div/PartRem[37][3] ,
         \u_div/PartRem[37][4] , \u_div/PartRem[37][5] ,
         \u_div/PartRem[38][0] , \u_div/PartRem[38][2] ,
         \u_div/PartRem[38][3] , \u_div/PartRem[38][4] ,
         \u_div/PartRem[38][5] , \u_div/PartRem[39][0] ,
         \u_div/PartRem[39][2] , \u_div/PartRem[39][3] ,
         \u_div/PartRem[39][4] , \u_div/PartRem[39][5] ,
         \u_div/PartRem[40][0] , \u_div/PartRem[40][2] ,
         \u_div/PartRem[40][3] , \u_div/PartRem[40][4] ,
         \u_div/PartRem[40][5] , \u_div/PartRem[41][0] ,
         \u_div/PartRem[41][2] , \u_div/PartRem[41][3] ,
         \u_div/PartRem[41][4] , \u_div/PartRem[41][5] ,
         \u_div/PartRem[42][0] , \u_div/PartRem[42][2] ,
         \u_div/PartRem[42][3] , \u_div/PartRem[42][4] ,
         \u_div/PartRem[42][5] , \u_div/PartRem[43][0] ,
         \u_div/PartRem[43][2] , \u_div/PartRem[43][3] ,
         \u_div/PartRem[43][4] , \u_div/PartRem[43][5] ,
         \u_div/PartRem[44][0] , \u_div/PartRem[44][2] ,
         \u_div/PartRem[44][3] , \u_div/PartRem[44][4] ,
         \u_div/PartRem[44][5] , \u_div/PartRem[45][0] ,
         \u_div/PartRem[45][2] , \u_div/PartRem[45][3] ,
         \u_div/PartRem[45][4] , \u_div/PartRem[45][5] ,
         \u_div/PartRem[46][0] , \u_div/PartRem[46][2] ,
         \u_div/PartRem[46][3] , \u_div/PartRem[46][4] ,
         \u_div/PartRem[46][5] , \u_div/PartRem[47][0] ,
         \u_div/PartRem[47][2] , \u_div/PartRem[47][3] ,
         \u_div/PartRem[47][4] , \u_div/PartRem[47][5] ,
         \u_div/PartRem[48][0] , \u_div/PartRem[48][2] ,
         \u_div/PartRem[48][3] , \u_div/PartRem[48][4] ,
         \u_div/PartRem[48][5] , \u_div/PartRem[49][0] ,
         \u_div/PartRem[49][2] , \u_div/PartRem[49][3] ,
         \u_div/PartRem[49][4] , \u_div/PartRem[49][5] ,
         \u_div/PartRem[50][0] , \u_div/PartRem[50][2] ,
         \u_div/PartRem[50][3] , \u_div/PartRem[50][4] ,
         \u_div/PartRem[50][5] , \u_div/PartRem[51][0] ,
         \u_div/PartRem[51][2] , \u_div/PartRem[51][3] ,
         \u_div/PartRem[51][4] , \u_div/PartRem[51][5] ,
         \u_div/PartRem[52][0] , \u_div/PartRem[52][2] ,
         \u_div/PartRem[52][3] , \u_div/PartRem[52][4] ,
         \u_div/PartRem[52][5] , \u_div/PartRem[53][0] ,
         \u_div/PartRem[53][2] , \u_div/PartRem[53][3] ,
         \u_div/PartRem[53][4] , \u_div/PartRem[53][5] ,
         \u_div/PartRem[54][0] , \u_div/PartRem[54][2] ,
         \u_div/PartRem[54][3] , \u_div/PartRem[54][4] ,
         \u_div/PartRem[54][5] , \u_div/PartRem[55][0] ,
         \u_div/PartRem[55][2] , \u_div/PartRem[55][3] ,
         \u_div/PartRem[55][4] , \u_div/PartRem[55][5] ,
         \u_div/PartRem[56][0] , \u_div/PartRem[56][2] ,
         \u_div/PartRem[56][3] , \u_div/PartRem[56][4] ,
         \u_div/PartRem[56][5] , \u_div/PartRem[57][0] ,
         \u_div/PartRem[57][2] , \u_div/PartRem[57][3] ,
         \u_div/PartRem[57][4] , \u_div/PartRem[57][5] ,
         \u_div/PartRem[58][0] , \u_div/PartRem[58][2] ,
         \u_div/PartRem[58][3] , \u_div/PartRem[58][4] ,
         \u_div/PartRem[58][5] , \u_div/PartRem[59][0] ,
         \u_div/PartRem[59][2] , \u_div/PartRem[59][3] ,
         \u_div/PartRem[59][4] , \u_div/PartRem[59][5] ,
         \u_div/PartRem[60][0] , \u_div/PartRem[61][0] ,
         \u_div/PartRem[62][0] , \u_div/PartRem[63][0] ,
         \u_div/PartRem[64][0] , \u_div/u_add_PartRem_2_1/n3 ,
         \u_div/u_add_PartRem_2_1/n2 , \u_div/u_add_PartRem_2_2/n3 ,
         \u_div/u_add_PartRem_2_2/n2 , \u_div/u_add_PartRem_2_3/n3 ,
         \u_div/u_add_PartRem_2_3/n2 , \u_div/u_add_PartRem_2_4/n3 ,
         \u_div/u_add_PartRem_2_4/n2 , \u_div/u_add_PartRem_2_5/n3 ,
         \u_div/u_add_PartRem_2_5/n2 , \u_div/u_add_PartRem_2_6/n3 ,
         \u_div/u_add_PartRem_2_6/n2 , \u_div/u_add_PartRem_2_7/n3 ,
         \u_div/u_add_PartRem_2_7/n2 , \u_div/u_add_PartRem_2_8/n3 ,
         \u_div/u_add_PartRem_2_8/n2 , \u_div/u_add_PartRem_2_9/n3 ,
         \u_div/u_add_PartRem_2_9/n2 , \u_div/u_add_PartRem_2_10/n3 ,
         \u_div/u_add_PartRem_2_10/n2 , \u_div/u_add_PartRem_2_11/n3 ,
         \u_div/u_add_PartRem_2_11/n2 , \u_div/u_add_PartRem_2_12/n3 ,
         \u_div/u_add_PartRem_2_12/n2 , \u_div/u_add_PartRem_2_13/n3 ,
         \u_div/u_add_PartRem_2_13/n2 , \u_div/u_add_PartRem_2_14/n3 ,
         \u_div/u_add_PartRem_2_14/n2 , \u_div/u_add_PartRem_2_15/n3 ,
         \u_div/u_add_PartRem_2_15/n2 , \u_div/u_add_PartRem_2_16/n3 ,
         \u_div/u_add_PartRem_2_16/n2 , \u_div/u_add_PartRem_2_17/n3 ,
         \u_div/u_add_PartRem_2_17/n2 , \u_div/u_add_PartRem_2_18/n3 ,
         \u_div/u_add_PartRem_2_18/n2 , \u_div/u_add_PartRem_2_19/n3 ,
         \u_div/u_add_PartRem_2_19/n2 , \u_div/u_add_PartRem_2_20/n3 ,
         \u_div/u_add_PartRem_2_20/n2 , \u_div/u_add_PartRem_2_21/n3 ,
         \u_div/u_add_PartRem_2_21/n2 , \u_div/u_add_PartRem_2_22/n3 ,
         \u_div/u_add_PartRem_2_22/n2 , \u_div/u_add_PartRem_2_23/n3 ,
         \u_div/u_add_PartRem_2_23/n2 , \u_div/u_add_PartRem_2_24/n3 ,
         \u_div/u_add_PartRem_2_24/n2 , \u_div/u_add_PartRem_2_25/n3 ,
         \u_div/u_add_PartRem_2_25/n2 , \u_div/u_add_PartRem_2_26/n3 ,
         \u_div/u_add_PartRem_2_26/n2 , \u_div/u_add_PartRem_2_27/n3 ,
         \u_div/u_add_PartRem_2_27/n2 , \u_div/u_add_PartRem_2_28/n3 ,
         \u_div/u_add_PartRem_2_28/n2 , \u_div/u_add_PartRem_2_29/n3 ,
         \u_div/u_add_PartRem_2_29/n2 , \u_div/u_add_PartRem_2_30/n3 ,
         \u_div/u_add_PartRem_2_30/n2 , \u_div/u_add_PartRem_2_31/n3 ,
         \u_div/u_add_PartRem_2_31/n2 , \u_div/u_add_PartRem_2_32/n3 ,
         \u_div/u_add_PartRem_2_32/n2 , \u_div/u_add_PartRem_2_33/n3 ,
         \u_div/u_add_PartRem_2_33/n2 , \u_div/u_add_PartRem_2_34/n3 ,
         \u_div/u_add_PartRem_2_34/n2 , \u_div/u_add_PartRem_2_35/n3 ,
         \u_div/u_add_PartRem_2_35/n2 , \u_div/u_add_PartRem_2_36/n3 ,
         \u_div/u_add_PartRem_2_36/n2 , \u_div/u_add_PartRem_2_37/n3 ,
         \u_div/u_add_PartRem_2_37/n2 , \u_div/u_add_PartRem_2_38/n3 ,
         \u_div/u_add_PartRem_2_38/n2 , \u_div/u_add_PartRem_2_39/n3 ,
         \u_div/u_add_PartRem_2_39/n2 , \u_div/u_add_PartRem_2_40/n3 ,
         \u_div/u_add_PartRem_2_40/n2 , \u_div/u_add_PartRem_2_41/n3 ,
         \u_div/u_add_PartRem_2_41/n2 , \u_div/u_add_PartRem_2_42/n3 ,
         \u_div/u_add_PartRem_2_42/n2 , \u_div/u_add_PartRem_2_43/n3 ,
         \u_div/u_add_PartRem_2_43/n2 , \u_div/u_add_PartRem_2_44/n3 ,
         \u_div/u_add_PartRem_2_44/n2 , \u_div/u_add_PartRem_2_45/n3 ,
         \u_div/u_add_PartRem_2_45/n2 , \u_div/u_add_PartRem_2_46/n3 ,
         \u_div/u_add_PartRem_2_46/n2 , \u_div/u_add_PartRem_2_47/n3 ,
         \u_div/u_add_PartRem_2_47/n2 , \u_div/u_add_PartRem_2_48/n3 ,
         \u_div/u_add_PartRem_2_48/n2 , \u_div/u_add_PartRem_2_49/n3 ,
         \u_div/u_add_PartRem_2_49/n2 , \u_div/u_add_PartRem_2_50/n3 ,
         \u_div/u_add_PartRem_2_50/n2 , \u_div/u_add_PartRem_2_51/n3 ,
         \u_div/u_add_PartRem_2_51/n2 , \u_div/u_add_PartRem_2_52/n3 ,
         \u_div/u_add_PartRem_2_52/n2 , \u_div/u_add_PartRem_2_53/n3 ,
         \u_div/u_add_PartRem_2_53/n2 , \u_div/u_add_PartRem_2_54/n3 ,
         \u_div/u_add_PartRem_2_54/n2 , \u_div/u_add_PartRem_2_55/n3 ,
         \u_div/u_add_PartRem_2_55/n2 , \u_div/u_add_PartRem_2_56/n3 ,
         \u_div/u_add_PartRem_2_56/n2 , \u_div/u_add_PartRem_2_57/n3 ,
         \u_div/u_add_PartRem_2_57/n2 , \u_div/u_add_PartRem_2_58/n3 ,
         \u_div/u_add_PartRem_2_58/n2 , n1, n2, n3, n4, n5, n6, n7, n8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign \u_div/QInv[63]  = a[63];

  GSIM_DW01_absval_3 \u_div/u_absval_AAbs  ( .A({n3, a[62:0]}), .ABSVAL({
        \u_div/PartRem[64][0] , \u_div/PartRem[63][0] , \u_div/PartRem[62][0] , 
        \u_div/PartRem[61][0] , \u_div/PartRem[60][0] , \u_div/PartRem[59][0] , 
        \u_div/PartRem[58][0] , \u_div/PartRem[57][0] , \u_div/PartRem[56][0] , 
        \u_div/PartRem[55][0] , \u_div/PartRem[54][0] , \u_div/PartRem[53][0] , 
        \u_div/PartRem[52][0] , \u_div/PartRem[51][0] , \u_div/PartRem[50][0] , 
        \u_div/PartRem[49][0] , \u_div/PartRem[48][0] , \u_div/PartRem[47][0] , 
        \u_div/PartRem[46][0] , \u_div/PartRem[45][0] , \u_div/PartRem[44][0] , 
        \u_div/PartRem[43][0] , \u_div/PartRem[42][0] , \u_div/PartRem[41][0] , 
        \u_div/PartRem[40][0] , \u_div/PartRem[39][0] , \u_div/PartRem[38][0] , 
        \u_div/PartRem[37][0] , \u_div/PartRem[36][0] , \u_div/PartRem[35][0] , 
        \u_div/PartRem[34][0] , \u_div/PartRem[33][0] , \u_div/PartRem[32][0] , 
        \u_div/PartRem[31][0] , \u_div/PartRem[30][0] , \u_div/PartRem[29][0] , 
        \u_div/PartRem[28][0] , \u_div/PartRem[27][0] , \u_div/PartRem[26][0] , 
        \u_div/PartRem[25][0] , \u_div/PartRem[24][0] , \u_div/PartRem[23][0] , 
        \u_div/PartRem[22][0] , \u_div/PartRem[21][0] , \u_div/PartRem[20][0] , 
        \u_div/PartRem[19][0] , \u_div/PartRem[18][0] , \u_div/PartRem[17][0] , 
        \u_div/PartRem[16][0] , \u_div/PartRem[15][0] , \u_div/PartRem[14][0] , 
        \u_div/PartRem[13][0] , \u_div/PartRem[12][0] , \u_div/PartRem[11][0] , 
        \u_div/PartRem[10][0] , \u_div/PartRem[9][0] , \u_div/PartRem[8][0] , 
        \u_div/PartRem[7][0] , \u_div/PartRem[6][0] , \u_div/PartRem[5][0] , 
        \u_div/PartRem[4][0] , \u_div/PartRem[3][0] , SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1}) );
  GSIM_DW_inc_3 \u_div/u_inc_QInc  ( .carry_in(n5), .a({n3, n3, n3, n4, 
        \u_div/QInv[59] , \u_div/QInv[58] , \u_div/QInv[57] , \u_div/QInv[56] , 
        \u_div/QInv[55] , \u_div/QInv[54] , \u_div/QInv[53] , \u_div/QInv[52] , 
        \u_div/QInv[51] , \u_div/QInv[50] , \u_div/QInv[49] , \u_div/QInv[48] , 
        \u_div/QInv[47] , \u_div/QInv[46] , \u_div/QInv[45] , \u_div/QInv[44] , 
        \u_div/QInv[43] , \u_div/QInv[42] , \u_div/QInv[41] , \u_div/QInv[40] , 
        \u_div/QInv[39] , \u_div/QInv[38] , \u_div/QInv[37] , \u_div/QInv[36] , 
        \u_div/QInv[35] , \u_div/QInv[34] , \u_div/QInv[33] , \u_div/QInv[32] , 
        \u_div/QInv[31] , \u_div/QInv[30] , \u_div/QInv[29] , \u_div/QInv[28] , 
        \u_div/QInv[27] , \u_div/QInv[26] , \u_div/QInv[25] , \u_div/QInv[24] , 
        \u_div/QInv[23] , \u_div/QInv[22] , \u_div/QInv[21] , \u_div/QInv[20] , 
        \u_div/QInv[19] , \u_div/QInv[18] , \u_div/QInv[17] , \u_div/QInv[16] , 
        \u_div/QInv[15] , \u_div/QInv[14] , \u_div/QInv[13] , \u_div/QInv[12] , 
        \u_div/QInv[11] , \u_div/QInv[10] , \u_div/QInv[9] , \u_div/QInv[8] , 
        \u_div/QInv[7] , \u_div/QInv[6] , \u_div/QInv[5] , \u_div/QInv[4] , 
        \u_div/QInv[3] , \u_div/QInv[2] , \u_div/QInv[1] , \u_div/QInv[0] }), 
        .sum(quotient) );
  ADDHXL \u_div/u_add_PartRem_2_2/U3  ( .A(\u_div/PartRem[3][4] ), .B(
        \u_div/u_add_PartRem_2_2/n3 ), .CO(\u_div/u_add_PartRem_2_2/n2 ), .S(
        \u_div/SumTmp[2][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_7/U3  ( .A(\u_div/PartRem[8][4] ), .B(
        \u_div/u_add_PartRem_2_7/n3 ), .CO(\u_div/u_add_PartRem_2_7/n2 ), .S(
        \u_div/SumTmp[7][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_12/U3  ( .A(\u_div/PartRem[13][4] ), .B(
        \u_div/u_add_PartRem_2_12/n3 ), .CO(\u_div/u_add_PartRem_2_12/n2 ), 
        .S(\u_div/SumTmp[12][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_17/U3  ( .A(\u_div/PartRem[18][4] ), .B(
        \u_div/u_add_PartRem_2_17/n3 ), .CO(\u_div/u_add_PartRem_2_17/n2 ), 
        .S(\u_div/SumTmp[17][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_22/U3  ( .A(\u_div/PartRem[23][4] ), .B(
        \u_div/u_add_PartRem_2_22/n3 ), .CO(\u_div/u_add_PartRem_2_22/n2 ), 
        .S(\u_div/SumTmp[22][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_27/U3  ( .A(\u_div/PartRem[28][4] ), .B(
        \u_div/u_add_PartRem_2_27/n3 ), .CO(\u_div/u_add_PartRem_2_27/n2 ), 
        .S(\u_div/SumTmp[27][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_32/U3  ( .A(\u_div/PartRem[33][4] ), .B(
        \u_div/u_add_PartRem_2_32/n3 ), .CO(\u_div/u_add_PartRem_2_32/n2 ), 
        .S(\u_div/SumTmp[32][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_37/U3  ( .A(\u_div/PartRem[38][4] ), .B(
        \u_div/u_add_PartRem_2_37/n3 ), .CO(\u_div/u_add_PartRem_2_37/n2 ), 
        .S(\u_div/SumTmp[37][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_42/U3  ( .A(\u_div/PartRem[43][4] ), .B(
        \u_div/u_add_PartRem_2_42/n3 ), .CO(\u_div/u_add_PartRem_2_42/n2 ), 
        .S(\u_div/SumTmp[42][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_47/U3  ( .A(\u_div/PartRem[48][4] ), .B(
        \u_div/u_add_PartRem_2_47/n3 ), .CO(\u_div/u_add_PartRem_2_47/n2 ), 
        .S(\u_div/SumTmp[47][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_52/U3  ( .A(\u_div/PartRem[53][4] ), .B(
        \u_div/u_add_PartRem_2_52/n3 ), .CO(\u_div/u_add_PartRem_2_52/n2 ), 
        .S(\u_div/SumTmp[52][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_53_1  ( .A(\u_div/SumTmp[53][1] ), .B(
        \u_div/SumTmp[53][1] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_48_1  ( .A(\u_div/SumTmp[48][1] ), .B(
        \u_div/SumTmp[48][1] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_43_1  ( .A(\u_div/SumTmp[43][1] ), .B(
        \u_div/SumTmp[43][1] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_38_1  ( .A(\u_div/SumTmp[38][1] ), .B(
        \u_div/SumTmp[38][1] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_33_1  ( .A(\u_div/SumTmp[33][1] ), .B(
        \u_div/SumTmp[33][1] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_28_1  ( .A(\u_div/SumTmp[28][1] ), .B(
        \u_div/SumTmp[28][1] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_23_1  ( .A(\u_div/SumTmp[23][1] ), .B(
        \u_div/SumTmp[23][1] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_0  ( .A(\u_div/PartRem[3][0] ), .B(
        \u_div/PartRem[3][0] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/SumTmp[1][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_0  ( .A(\u_div/PartRem[22][0] ), .B(
        \u_div/PartRem[22][0] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/SumTmp[20][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_20_1  ( .A(\u_div/SumTmp[20][1] ), .B(
        \u_div/SumTmp[20][1] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_0  ( .A(\u_div/PartRem[6][0] ), .B(
        \u_div/PartRem[6][0] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/SumTmp[4][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_0  ( .A(\u_div/PartRem[7][0] ), .B(
        \u_div/PartRem[7][0] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/SumTmp[5][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_0  ( .A(\u_div/PartRem[12][0] ), .B(
        \u_div/PartRem[12][0] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/SumTmp[10][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_0  ( .A(\u_div/PartRem[13][0] ), .B(
        \u_div/PartRem[13][0] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/SumTmp[11][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_0  ( .A(\u_div/PartRem[16][0] ), .B(
        \u_div/PartRem[16][0] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/SumTmp[14][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_0  ( .A(\u_div/PartRem[17][0] ), .B(
        \u_div/PartRem[17][0] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/SumTmp[15][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_0  ( .A(\u_div/PartRem[19][0] ), .B(
        \u_div/PartRem[19][0] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/SumTmp[17][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_0  ( .A(\u_div/PartRem[23][0] ), .B(
        \u_div/PartRem[23][0] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/SumTmp[21][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_0  ( .A(\u_div/PartRem[26][0] ), .B(
        \u_div/PartRem[26][0] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/SumTmp[24][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_0  ( .A(\u_div/PartRem[27][0] ), .B(
        \u_div/PartRem[27][0] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/SumTmp[25][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_0  ( .A(\u_div/PartRem[28][0] ), .B(
        \u_div/PartRem[28][0] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/SumTmp[26][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_0  ( .A(\u_div/PartRem[31][0] ), .B(
        \u_div/PartRem[31][0] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/SumTmp[29][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_0  ( .A(\u_div/PartRem[32][0] ), .B(
        \u_div/PartRem[32][0] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/SumTmp[30][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_0  ( .A(\u_div/PartRem[33][0] ), .B(
        \u_div/PartRem[33][0] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/SumTmp[31][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_0  ( .A(\u_div/PartRem[36][0] ), .B(
        \u_div/PartRem[36][0] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/SumTmp[34][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_0  ( .A(\u_div/PartRem[37][0] ), .B(
        \u_div/PartRem[37][0] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/SumTmp[35][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_0  ( .A(\u_div/PartRem[38][0] ), .B(
        \u_div/PartRem[38][0] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/SumTmp[36][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_0  ( .A(\u_div/PartRem[41][0] ), .B(
        \u_div/PartRem[41][0] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/SumTmp[39][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_0  ( .A(\u_div/PartRem[42][0] ), .B(
        \u_div/PartRem[42][0] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/SumTmp[40][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_0  ( .A(\u_div/PartRem[43][0] ), .B(
        \u_div/PartRem[43][0] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/SumTmp[41][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_0  ( .A(\u_div/PartRem[46][0] ), .B(
        \u_div/PartRem[46][0] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/SumTmp[44][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_0  ( .A(\u_div/PartRem[47][0] ), .B(
        \u_div/PartRem[47][0] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/SumTmp[45][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_0  ( .A(\u_div/PartRem[48][0] ), .B(
        \u_div/PartRem[48][0] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/SumTmp[46][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_0  ( .A(\u_div/PartRem[51][0] ), .B(
        \u_div/PartRem[51][0] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/SumTmp[49][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_0  ( .A(\u_div/PartRem[52][0] ), .B(
        \u_div/PartRem[52][0] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/SumTmp[50][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_0  ( .A(\u_div/PartRem[53][0] ), .B(
        \u_div/PartRem[53][0] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/SumTmp[51][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_0  ( .A(\u_div/PartRem[56][0] ), .B(
        \u_div/PartRem[56][0] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/SumTmp[54][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_0  ( .A(\u_div/PartRem[57][0] ), .B(
        \u_div/PartRem[57][0] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/SumTmp[55][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_0  ( .A(\u_div/PartRem[59][0] ), .B(
        \u_div/PartRem[59][0] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/SumTmp[57][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_0  ( .A(\u_div/PartRem[60][0] ), .B(
        \u_div/PartRem[60][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/SumTmp[58][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_9_0  ( .A(\u_div/PartRem[10][0] ), .B(
        \u_div/PartRem[10][0] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/SumTmp[8][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_0  ( .A(\u_div/PartRem[15][0] ), .B(
        \u_div/PartRem[15][0] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/SumTmp[13][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_0  ( .A(\u_div/PartRem[20][0] ), .B(
        \u_div/PartRem[20][0] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/SumTmp[18][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_0  ( .A(\u_div/PartRem[4][0] ), .B(
        \u_div/PartRem[4][0] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/SumTmp[2][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_0  ( .A(\u_div/PartRem[5][0] ), .B(
        \u_div/PartRem[5][0] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/SumTmp[3][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_59_1  ( .A(\u_div/PartRem[61][0] ), .B(
        \u_div/PartRem[61][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_0  ( .A(\u_div/PartRem[8][0] ), .B(
        \u_div/PartRem[8][0] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/SumTmp[6][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_0  ( .A(\u_div/PartRem[11][0] ), .B(
        \u_div/PartRem[11][0] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/SumTmp[9][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_0  ( .A(\u_div/PartRem[14][0] ), .B(
        \u_div/PartRem[14][0] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/SumTmp[12][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_0  ( .A(\u_div/PartRem[18][0] ), .B(
        \u_div/PartRem[18][0] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/SumTmp[16][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_0  ( .A(\u_div/PartRem[58][0] ), .B(
        \u_div/PartRem[58][0] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/SumTmp[56][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_0  ( .A(\u_div/PartRem[25][0] ), .B(
        \u_div/PartRem[25][0] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/SumTmp[23][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_0  ( .A(\u_div/PartRem[30][0] ), .B(
        \u_div/PartRem[30][0] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/SumTmp[28][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_0  ( .A(\u_div/PartRem[35][0] ), .B(
        \u_div/PartRem[35][0] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/SumTmp[33][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_0  ( .A(\u_div/PartRem[40][0] ), .B(
        \u_div/PartRem[40][0] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/SumTmp[38][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_0  ( .A(\u_div/PartRem[45][0] ), .B(
        \u_div/PartRem[45][0] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/SumTmp[43][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_0  ( .A(\u_div/PartRem[50][0] ), .B(
        \u_div/PartRem[50][0] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/SumTmp[48][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_0  ( .A(\u_div/PartRem[55][0] ), .B(
        \u_div/PartRem[55][0] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/SumTmp[53][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_3  ( .A(\u_div/PartRem[4][3] ), .B(
        \u_div/SumTmp[3][3] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_3  ( .A(\u_div/PartRem[6][3] ), .B(
        \u_div/SumTmp[5][3] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_3  ( .A(\u_div/PartRem[8][3] ), .B(
        \u_div/SumTmp[7][3] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_8_3  ( .A(\u_div/PartRem[9][3] ), .B(
        \u_div/SumTmp[8][3] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_3  ( .A(\u_div/PartRem[11][3] ), .B(
        \u_div/SumTmp[10][3] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_3  ( .A(\u_div/PartRem[12][3] ), .B(
        \u_div/SumTmp[11][3] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_3  ( .A(\u_div/PartRem[14][3] ), .B(
        \u_div/SumTmp[13][3] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_3  ( .A(\u_div/PartRem[15][3] ), .B(
        \u_div/SumTmp[14][3] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_3  ( .A(\u_div/PartRem[16][3] ), .B(
        \u_div/SumTmp[15][3] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_3  ( .A(\u_div/PartRem[18][3] ), .B(
        \u_div/SumTmp[17][3] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_3  ( .A(\u_div/PartRem[19][3] ), .B(
        \u_div/SumTmp[18][3] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_3  ( .A(\u_div/PartRem[22][3] ), .B(
        \u_div/SumTmp[21][3] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_3  ( .A(\u_div/PartRem[23][3] ), .B(
        \u_div/SumTmp[22][3] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_3  ( .A(\u_div/PartRem[25][3] ), .B(
        \u_div/SumTmp[24][3] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_3  ( .A(\u_div/PartRem[26][3] ), .B(
        \u_div/SumTmp[25][3] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_3  ( .A(\u_div/PartRem[28][3] ), .B(
        \u_div/SumTmp[27][3] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_3  ( .A(\u_div/PartRem[30][3] ), .B(
        \u_div/SumTmp[29][3] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_3  ( .A(\u_div/PartRem[31][3] ), .B(
        \u_div/SumTmp[30][3] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_3  ( .A(\u_div/PartRem[33][3] ), .B(
        \u_div/SumTmp[32][3] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_3  ( .A(\u_div/PartRem[35][3] ), .B(
        \u_div/SumTmp[34][3] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_3  ( .A(\u_div/PartRem[36][3] ), .B(
        \u_div/SumTmp[35][3] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_3  ( .A(\u_div/PartRem[38][3] ), .B(
        \u_div/SumTmp[37][3] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_3  ( .A(\u_div/PartRem[40][3] ), .B(
        \u_div/SumTmp[39][3] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_3  ( .A(\u_div/PartRem[41][3] ), .B(
        \u_div/SumTmp[40][3] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_3  ( .A(\u_div/PartRem[43][3] ), .B(
        \u_div/SumTmp[42][3] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_3  ( .A(\u_div/PartRem[45][3] ), .B(
        \u_div/SumTmp[44][3] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_3  ( .A(\u_div/PartRem[46][3] ), .B(
        \u_div/SumTmp[45][3] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_3  ( .A(\u_div/PartRem[48][3] ), .B(
        \u_div/SumTmp[47][3] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_3  ( .A(\u_div/PartRem[50][3] ), .B(
        \u_div/SumTmp[49][3] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_3  ( .A(\u_div/PartRem[51][3] ), .B(
        \u_div/SumTmp[50][3] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_3  ( .A(\u_div/PartRem[53][3] ), .B(
        \u_div/SumTmp[52][3] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_3  ( .A(\u_div/PartRem[55][3] ), .B(
        \u_div/SumTmp[54][3] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_3  ( .A(\u_div/PartRem[56][3] ), .B(
        \u_div/SumTmp[55][3] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_3  ( .A(\u_div/PartRem[58][3] ), .B(
        \u_div/SumTmp[57][3] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_3  ( .A(\u_div/PartRem[59][3] ), .B(
        \u_div/SumTmp[58][3] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_3  ( .A(\u_div/PartRem[5][3] ), .B(
        \u_div/SumTmp[4][3] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_3  ( .A(\u_div/PartRem[27][3] ), .B(
        \u_div/SumTmp[26][3] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_3  ( .A(\u_div/PartRem[32][3] ), .B(
        \u_div/SumTmp[31][3] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_3  ( .A(\u_div/PartRem[37][3] ), .B(
        \u_div/SumTmp[36][3] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_3  ( .A(\u_div/PartRem[42][3] ), .B(
        \u_div/SumTmp[41][3] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_3  ( .A(\u_div/PartRem[47][3] ), .B(
        \u_div/SumTmp[46][3] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_3  ( .A(\u_div/PartRem[52][3] ), .B(
        \u_div/SumTmp[51][3] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_3  ( .A(\u_div/PartRem[63][0] ), .B(
        \u_div/SumTmp[59][3] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_3  ( .A(\u_div/PartRem[3][3] ), .B(
        \u_div/SumTmp[2][3] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_3  ( .A(\u_div/PartRem[7][3] ), .B(
        \u_div/SumTmp[6][3] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_9_3  ( .A(\u_div/PartRem[10][3] ), .B(
        \u_div/SumTmp[9][3] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_3  ( .A(\u_div/PartRem[13][3] ), .B(
        \u_div/SumTmp[12][3] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_3  ( .A(\u_div/PartRem[17][3] ), .B(
        \u_div/SumTmp[16][3] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_3  ( .A(\u_div/PartRem[20][3] ), .B(
        \u_div/SumTmp[19][3] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_3  ( .A(\u_div/PartRem[57][3] ), .B(
        \u_div/SumTmp[56][3] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_4  ( .A(\u_div/PartRem[64][0] ), .B(
        \u_div/SumTmp[59][4] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_3_1  ( .A(\u_div/SumTmp[3][1] ), .B(
        \u_div/SumTmp[3][1] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_4_1  ( .A(\u_div/SumTmp[4][1] ), .B(
        \u_div/SumTmp[4][1] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_5_1  ( .A(\u_div/SumTmp[5][1] ), .B(
        \u_div/SumTmp[5][1] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_6_1  ( .A(\u_div/SumTmp[6][1] ), .B(
        \u_div/SumTmp[6][1] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_7_1  ( .A(\u_div/SumTmp[7][1] ), .B(
        \u_div/SumTmp[7][1] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_9_1  ( .A(\u_div/SumTmp[9][1] ), .B(
        \u_div/SumTmp[9][1] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_10_1  ( .A(\u_div/SumTmp[10][1] ), .B(
        \u_div/SumTmp[10][1] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_11_1  ( .A(\u_div/SumTmp[11][1] ), .B(
        \u_div/SumTmp[11][1] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_12_1  ( .A(\u_div/SumTmp[12][1] ), .B(
        \u_div/SumTmp[12][1] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_13_1  ( .A(\u_div/SumTmp[13][1] ), .B(
        \u_div/SumTmp[13][1] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_14_1  ( .A(\u_div/SumTmp[14][1] ), .B(
        \u_div/SumTmp[14][1] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_15_1  ( .A(\u_div/SumTmp[15][1] ), .B(
        \u_div/SumTmp[15][1] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_16_1  ( .A(\u_div/SumTmp[16][1] ), .B(
        \u_div/SumTmp[16][1] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_17_1  ( .A(\u_div/SumTmp[17][1] ), .B(
        \u_div/SumTmp[17][1] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_18_1  ( .A(\u_div/SumTmp[18][1] ), .B(
        \u_div/SumTmp[18][1] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_19_1  ( .A(\u_div/SumTmp[19][1] ), .B(
        \u_div/SumTmp[19][1] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_0  ( .A(\u_div/PartRem[21][0] ), .B(
        \u_div/PartRem[21][0] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/SumTmp[19][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_22_1  ( .A(\u_div/SumTmp[22][1] ), .B(
        \u_div/SumTmp[22][1] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_0  ( .A(\u_div/PartRem[24][0] ), .B(
        \u_div/PartRem[24][0] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/SumTmp[22][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_21_1  ( .A(\u_div/SumTmp[21][1] ), .B(
        \u_div/SumTmp[21][1] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_25_1  ( .A(\u_div/SumTmp[25][1] ), .B(
        \u_div/SumTmp[25][1] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_26_1  ( .A(\u_div/SumTmp[26][1] ), .B(
        \u_div/SumTmp[26][1] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_24_1  ( .A(\u_div/SumTmp[24][1] ), .B(
        \u_div/SumTmp[24][1] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_27_1  ( .A(\u_div/SumTmp[27][1] ), .B(
        \u_div/SumTmp[27][1] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_0  ( .A(\u_div/PartRem[29][0] ), .B(
        \u_div/PartRem[29][0] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/SumTmp[27][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_29_1  ( .A(\u_div/SumTmp[29][1] ), .B(
        \u_div/SumTmp[29][1] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_30_1  ( .A(\u_div/SumTmp[30][1] ), .B(
        \u_div/SumTmp[30][1] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_31_1  ( .A(\u_div/SumTmp[31][1] ), .B(
        \u_div/SumTmp[31][1] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_32_1  ( .A(\u_div/SumTmp[32][1] ), .B(
        \u_div/SumTmp[32][1] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_0  ( .A(\u_div/PartRem[34][0] ), .B(
        \u_div/PartRem[34][0] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/SumTmp[32][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_34_1  ( .A(\u_div/SumTmp[34][1] ), .B(
        \u_div/SumTmp[34][1] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_35_1  ( .A(\u_div/SumTmp[35][1] ), .B(
        \u_div/SumTmp[35][1] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_36_1  ( .A(\u_div/SumTmp[36][1] ), .B(
        \u_div/SumTmp[36][1] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_37_1  ( .A(\u_div/SumTmp[37][1] ), .B(
        \u_div/SumTmp[37][1] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_0  ( .A(\u_div/PartRem[39][0] ), .B(
        \u_div/PartRem[39][0] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/SumTmp[37][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_39_1  ( .A(\u_div/SumTmp[39][1] ), .B(
        \u_div/SumTmp[39][1] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_40_1  ( .A(\u_div/SumTmp[40][1] ), .B(
        \u_div/SumTmp[40][1] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_41_1  ( .A(\u_div/SumTmp[41][1] ), .B(
        \u_div/SumTmp[41][1] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_42_1  ( .A(\u_div/SumTmp[42][1] ), .B(
        \u_div/SumTmp[42][1] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_0  ( .A(\u_div/PartRem[44][0] ), .B(
        \u_div/PartRem[44][0] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/SumTmp[42][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_44_1  ( .A(\u_div/SumTmp[44][1] ), .B(
        \u_div/SumTmp[44][1] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_45_1  ( .A(\u_div/SumTmp[45][1] ), .B(
        \u_div/SumTmp[45][1] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_46_1  ( .A(\u_div/SumTmp[46][1] ), .B(
        \u_div/SumTmp[46][1] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_47_1  ( .A(\u_div/SumTmp[47][1] ), .B(
        \u_div/SumTmp[47][1] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_0  ( .A(\u_div/PartRem[49][0] ), .B(
        \u_div/PartRem[49][0] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/SumTmp[47][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_49_1  ( .A(\u_div/SumTmp[49][1] ), .B(
        \u_div/SumTmp[49][1] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_51_1  ( .A(\u_div/SumTmp[51][1] ), .B(
        \u_div/SumTmp[51][1] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_50_1  ( .A(\u_div/SumTmp[50][1] ), .B(
        \u_div/SumTmp[50][1] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_52_1  ( .A(\u_div/SumTmp[52][1] ), .B(
        \u_div/SumTmp[52][1] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_0  ( .A(\u_div/PartRem[54][0] ), .B(
        \u_div/PartRem[54][0] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/SumTmp[52][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_54_1  ( .A(\u_div/SumTmp[54][1] ), .B(
        \u_div/SumTmp[54][1] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_55_1  ( .A(\u_div/SumTmp[55][1] ), .B(
        \u_div/SumTmp[55][1] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_56_1  ( .A(\u_div/SumTmp[56][1] ), .B(
        \u_div/SumTmp[56][1] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_57_1  ( .A(\u_div/SumTmp[57][1] ), .B(
        \u_div/SumTmp[57][1] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_58_1  ( .A(\u_div/SumTmp[58][1] ), .B(
        \u_div/SumTmp[58][1] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_3  ( .A(\u_div/PartRem[21][3] ), .B(
        \u_div/SumTmp[20][3] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_3  ( .A(\u_div/PartRem[24][3] ), .B(
        \u_div/SumTmp[23][3] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_3  ( .A(\u_div/PartRem[29][3] ), .B(
        \u_div/SumTmp[28][3] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_3  ( .A(\u_div/PartRem[34][3] ), .B(
        \u_div/SumTmp[33][3] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_3  ( .A(\u_div/PartRem[39][3] ), .B(
        \u_div/SumTmp[38][3] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_3  ( .A(\u_div/PartRem[44][3] ), .B(
        \u_div/SumTmp[43][3] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_3  ( .A(\u_div/PartRem[49][3] ), .B(
        \u_div/SumTmp[48][3] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_3  ( .A(\u_div/PartRem[54][3] ), .B(
        \u_div/SumTmp[53][3] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_1_3  ( .A(\u_div/PartRem[2][3] ), .B(
        \u_div/SumTmp[1][3] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][4] ) );
  MX2X1 \u_div/u_mx_PartRem_1_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/SumTmp[1][2] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][3] ) );
  MX2XL \u_div/u_mx_PartRem_1_1_4  ( .A(\u_div/PartRem[2][4] ), .B(
        \u_div/SumTmp[1][4] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_4  ( .A(\u_div/PartRem[22][4] ), .B(
        \u_div/SumTmp[21][4] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_4  ( .A(\u_div/PartRem[25][4] ), .B(
        \u_div/SumTmp[24][4] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_4  ( .A(\u_div/PartRem[30][4] ), .B(
        \u_div/SumTmp[29][4] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_4  ( .A(\u_div/PartRem[35][4] ), .B(
        \u_div/SumTmp[34][4] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_4  ( .A(\u_div/PartRem[40][4] ), .B(
        \u_div/SumTmp[39][4] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_4  ( .A(\u_div/PartRem[50][4] ), .B(
        \u_div/SumTmp[49][4] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_4  ( .A(\u_div/PartRem[45][4] ), .B(
        \u_div/SumTmp[44][4] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_4  ( .A(\u_div/PartRem[55][4] ), .B(
        \u_div/SumTmp[54][4] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_4  ( .A(\u_div/PartRem[3][4] ), .B(
        \u_div/SumTmp[2][4] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_4  ( .A(\u_div/PartRem[4][4] ), .B(
        \u_div/SumTmp[3][4] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_4  ( .A(\u_div/PartRem[5][4] ), .B(
        \u_div/SumTmp[4][4] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_4  ( .A(\u_div/PartRem[6][4] ), .B(
        \u_div/SumTmp[5][4] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_4  ( .A(\u_div/PartRem[7][4] ), .B(
        \u_div/SumTmp[6][4] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_4  ( .A(\u_div/PartRem[8][4] ), .B(
        \u_div/SumTmp[7][4] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_9_4  ( .A(\u_div/PartRem[10][4] ), .B(
        \u_div/SumTmp[9][4] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_4  ( .A(\u_div/PartRem[11][4] ), .B(
        \u_div/SumTmp[10][4] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_4  ( .A(\u_div/PartRem[12][4] ), .B(
        \u_div/SumTmp[11][4] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_4  ( .A(\u_div/PartRem[13][4] ), .B(
        \u_div/SumTmp[12][4] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_4  ( .A(\u_div/PartRem[14][4] ), .B(
        \u_div/SumTmp[13][4] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_4  ( .A(\u_div/PartRem[15][4] ), .B(
        \u_div/SumTmp[14][4] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_4  ( .A(\u_div/PartRem[16][4] ), .B(
        \u_div/SumTmp[15][4] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_4  ( .A(\u_div/PartRem[17][4] ), .B(
        \u_div/SumTmp[16][4] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_4  ( .A(\u_div/PartRem[18][4] ), .B(
        \u_div/SumTmp[17][4] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_4  ( .A(\u_div/PartRem[19][4] ), .B(
        \u_div/SumTmp[18][4] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_4  ( .A(\u_div/PartRem[20][4] ), .B(
        \u_div/SumTmp[19][4] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_4  ( .A(\u_div/PartRem[21][4] ), .B(
        \u_div/SumTmp[20][4] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_4  ( .A(\u_div/PartRem[23][4] ), .B(
        \u_div/SumTmp[22][4] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_4  ( .A(\u_div/PartRem[26][4] ), .B(
        \u_div/SumTmp[25][4] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_4  ( .A(\u_div/PartRem[24][4] ), .B(
        \u_div/SumTmp[23][4] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_4  ( .A(\u_div/PartRem[29][4] ), .B(
        \u_div/SumTmp[28][4] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_4  ( .A(\u_div/PartRem[27][4] ), .B(
        \u_div/SumTmp[26][4] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_4  ( .A(\u_div/PartRem[28][4] ), .B(
        \u_div/SumTmp[27][4] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_4  ( .A(\u_div/PartRem[31][4] ), .B(
        \u_div/SumTmp[30][4] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_4  ( .A(\u_div/PartRem[34][4] ), .B(
        \u_div/SumTmp[33][4] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_4  ( .A(\u_div/PartRem[32][4] ), .B(
        \u_div/SumTmp[31][4] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_4  ( .A(\u_div/PartRem[33][4] ), .B(
        \u_div/SumTmp[32][4] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_4  ( .A(\u_div/PartRem[36][4] ), .B(
        \u_div/SumTmp[35][4] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_4  ( .A(\u_div/PartRem[37][4] ), .B(
        \u_div/SumTmp[36][4] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_4  ( .A(\u_div/PartRem[39][4] ), .B(
        \u_div/SumTmp[38][4] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_4  ( .A(\u_div/PartRem[38][4] ), .B(
        \u_div/SumTmp[37][4] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_4  ( .A(\u_div/PartRem[41][4] ), .B(
        \u_div/SumTmp[40][4] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_4  ( .A(\u_div/PartRem[44][4] ), .B(
        \u_div/SumTmp[43][4] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_4  ( .A(\u_div/PartRem[42][4] ), .B(
        \u_div/SumTmp[41][4] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_4  ( .A(\u_div/PartRem[43][4] ), .B(
        \u_div/SumTmp[42][4] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_4  ( .A(\u_div/PartRem[47][4] ), .B(
        \u_div/SumTmp[46][4] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_4  ( .A(\u_div/PartRem[46][4] ), .B(
        \u_div/SumTmp[45][4] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_4  ( .A(\u_div/PartRem[52][4] ), .B(
        \u_div/SumTmp[51][4] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_4  ( .A(\u_div/PartRem[48][4] ), .B(
        \u_div/SumTmp[47][4] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_4  ( .A(\u_div/PartRem[49][4] ), .B(
        \u_div/SumTmp[48][4] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_4  ( .A(\u_div/PartRem[51][4] ), .B(
        \u_div/SumTmp[50][4] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_4  ( .A(\u_div/PartRem[53][4] ), .B(
        \u_div/SumTmp[52][4] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_4  ( .A(\u_div/PartRem[54][4] ), .B(
        \u_div/SumTmp[53][4] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_4  ( .A(\u_div/PartRem[58][4] ), .B(
        \u_div/SumTmp[57][4] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_4  ( .A(\u_div/PartRem[56][4] ), .B(
        \u_div/SumTmp[55][4] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_4  ( .A(\u_div/PartRem[57][4] ), .B(
        \u_div/SumTmp[56][4] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_4  ( .A(\u_div/PartRem[59][4] ), .B(
        \u_div/SumTmp[58][4] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_8_4  ( .A(\u_div/PartRem[9][4] ), .B(
        \u_div/SumTmp[8][4] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][5] ) );
  CLKMX2X6 \u_div/u_mx_PartRem_1_8_1  ( .A(\u_div/SumTmp[8][1] ), .B(
        \u_div/SumTmp[8][1] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_8_0  ( .A(\u_div/PartRem[9][0] ), .B(
        \u_div/PartRem[9][0] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/SumTmp[7][1] ) );
  MX2X6 \u_div/u_mx_PartRem_1_2_1  ( .A(\u_div/SumTmp[2][1] ), .B(
        \u_div/SumTmp[2][1] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][2] ) );
  OR2X2 U1 ( .A(\u_div/PartRem[8][5] ), .B(\u_div/u_add_PartRem_2_7/n2 ), .Y(
        \u_div/CryTmp[7][6] ) );
  XOR2XL U2 ( .A(\u_div/CryTmp[2][6] ), .B(n3), .Y(\u_div/QInv[2] ) );
  MXI2X4 U3 ( .A(\u_div/SumTmp[2][2] ), .B(\u_div/PartRem[3][2] ), .S0(
        \u_div/CryTmp[2][6] ), .Y(\u_div/PartRem[2][3] ) );
  OR2X6 U4 ( .A(\u_div/PartRem[3][5] ), .B(\u_div/u_add_PartRem_2_2/n2 ), .Y(
        \u_div/CryTmp[2][6] ) );
  OR2X8 U5 ( .A(\u_div/PartRem[52][5] ), .B(\u_div/u_add_PartRem_2_51/n2 ), 
        .Y(\u_div/CryTmp[51][6] ) );
  ADDHX2 U6 ( .A(\u_div/PartRem[52][4] ), .B(\u_div/u_add_PartRem_2_51/n3 ), 
        .CO(\u_div/u_add_PartRem_2_51/n2 ), .S(\u_div/SumTmp[51][4] ) );
  OR2X8 U7 ( .A(\u_div/PartRem[14][5] ), .B(\u_div/u_add_PartRem_2_13/n2 ), 
        .Y(\u_div/CryTmp[13][6] ) );
  ADDHX2 U8 ( .A(\u_div/PartRem[14][4] ), .B(\u_div/u_add_PartRem_2_13/n3 ), 
        .CO(\u_div/u_add_PartRem_2_13/n2 ), .S(\u_div/SumTmp[13][4] ) );
  OR2X8 U9 ( .A(\u_div/PartRem[5][5] ), .B(\u_div/u_add_PartRem_2_4/n2 ), .Y(
        \u_div/CryTmp[4][6] ) );
  ADDHX2 U10 ( .A(\u_div/PartRem[5][4] ), .B(\u_div/u_add_PartRem_2_4/n3 ), 
        .CO(\u_div/u_add_PartRem_2_4/n2 ), .S(\u_div/SumTmp[4][4] ) );
  MXI2X1 U11 ( .A(\u_div/SumTmp[31][2] ), .B(\u_div/PartRem[32][2] ), .S0(
        \u_div/CryTmp[31][6] ), .Y(\u_div/PartRem[31][3] ) );
  MXI2X1 U12 ( .A(\u_div/SumTmp[41][2] ), .B(\u_div/PartRem[42][2] ), .S0(
        \u_div/CryTmp[41][6] ), .Y(\u_div/PartRem[41][3] ) );
  OR2X1 U13 ( .A(\u_div/PartRem[12][2] ), .B(\u_div/PartRem[12][3] ), .Y(
        \u_div/u_add_PartRem_2_11/n3 ) );
  OR2X1 U14 ( .A(\u_div/PartRem[15][2] ), .B(\u_div/PartRem[15][3] ), .Y(
        \u_div/u_add_PartRem_2_14/n3 ) );
  OR2X1 U15 ( .A(\u_div/PartRem[16][2] ), .B(\u_div/PartRem[16][3] ), .Y(
        \u_div/u_add_PartRem_2_15/n3 ) );
  OR2X1 U16 ( .A(\u_div/PartRem[17][2] ), .B(\u_div/PartRem[17][3] ), .Y(
        \u_div/u_add_PartRem_2_16/n3 ) );
  MXI2X1 U17 ( .A(\u_div/SumTmp[3][2] ), .B(\u_div/PartRem[4][2] ), .S0(
        \u_div/CryTmp[3][6] ), .Y(\u_div/PartRem[3][3] ) );
  OR2X1 U18 ( .A(\u_div/PartRem[7][2] ), .B(\u_div/PartRem[7][3] ), .Y(
        \u_div/u_add_PartRem_2_6/n3 ) );
  OR2X1 U19 ( .A(\u_div/PartRem[11][2] ), .B(\u_div/PartRem[11][3] ), .Y(
        \u_div/u_add_PartRem_2_10/n3 ) );
  OR2X1 U20 ( .A(\u_div/PartRem[6][2] ), .B(\u_div/PartRem[6][3] ), .Y(
        \u_div/u_add_PartRem_2_5/n3 ) );
  OR2X1 U21 ( .A(\u_div/PartRem[5][2] ), .B(\u_div/PartRem[5][3] ), .Y(
        \u_div/u_add_PartRem_2_4/n3 ) );
  OR2X1 U22 ( .A(\u_div/PartRem[25][2] ), .B(\u_div/PartRem[25][3] ), .Y(
        \u_div/u_add_PartRem_2_24/n3 ) );
  OR2X1 U23 ( .A(\u_div/PartRem[29][2] ), .B(\u_div/PartRem[29][3] ), .Y(
        \u_div/u_add_PartRem_2_28/n3 ) );
  OR2X1 U24 ( .A(\u_div/PartRem[32][2] ), .B(\u_div/PartRem[32][3] ), .Y(
        \u_div/u_add_PartRem_2_31/n3 ) );
  OR2X1 U25 ( .A(\u_div/PartRem[34][2] ), .B(\u_div/PartRem[34][3] ), .Y(
        \u_div/u_add_PartRem_2_33/n3 ) );
  OR2X1 U26 ( .A(\u_div/PartRem[35][2] ), .B(\u_div/PartRem[35][3] ), .Y(
        \u_div/u_add_PartRem_2_34/n3 ) );
  OR2X1 U27 ( .A(\u_div/PartRem[39][2] ), .B(\u_div/PartRem[39][3] ), .Y(
        \u_div/u_add_PartRem_2_38/n3 ) );
  OR2X1 U28 ( .A(\u_div/PartRem[42][2] ), .B(\u_div/PartRem[42][3] ), .Y(
        \u_div/u_add_PartRem_2_41/n3 ) );
  OR2X1 U29 ( .A(\u_div/PartRem[44][2] ), .B(\u_div/PartRem[44][3] ), .Y(
        \u_div/u_add_PartRem_2_43/n3 ) );
  OR2X1 U30 ( .A(\u_div/PartRem[45][2] ), .B(\u_div/PartRem[45][3] ), .Y(
        \u_div/u_add_PartRem_2_44/n3 ) );
  OR2X1 U31 ( .A(\u_div/PartRem[50][2] ), .B(\u_div/PartRem[50][3] ), .Y(
        \u_div/u_add_PartRem_2_49/n3 ) );
  OR2X1 U32 ( .A(\u_div/PartRem[49][2] ), .B(\u_div/PartRem[49][3] ), .Y(
        \u_div/u_add_PartRem_2_48/n3 ) );
  OR2X1 U33 ( .A(\u_div/PartRem[52][2] ), .B(\u_div/PartRem[52][3] ), .Y(
        \u_div/u_add_PartRem_2_51/n3 ) );
  OR2X1 U34 ( .A(\u_div/PartRem[54][2] ), .B(\u_div/PartRem[54][3] ), .Y(
        \u_div/u_add_PartRem_2_53/n3 ) );
  OR2X1 U35 ( .A(\u_div/PartRem[55][2] ), .B(\u_div/PartRem[55][3] ), .Y(
        \u_div/u_add_PartRem_2_54/n3 ) );
  OR2X1 U36 ( .A(\u_div/PartRem[57][2] ), .B(\u_div/PartRem[57][3] ), .Y(
        \u_div/u_add_PartRem_2_56/n3 ) );
  OR2X1 U37 ( .A(\u_div/PartRem[58][2] ), .B(\u_div/PartRem[58][3] ), .Y(
        \u_div/u_add_PartRem_2_57/n3 ) );
  NOR2X1 U38 ( .A(\u_div/PartRem[63][0] ), .B(\u_div/PartRem[62][0] ), .Y(n8)
         );
  OR2X2 U39 ( .A(\u_div/PartRem[19][5] ), .B(\u_div/u_add_PartRem_2_18/n2 ), 
        .Y(\u_div/CryTmp[18][6] ) );
  OR2X2 U40 ( .A(\u_div/PartRem[21][5] ), .B(\u_div/u_add_PartRem_2_20/n2 ), 
        .Y(\u_div/CryTmp[20][6] ) );
  OR2X2 U41 ( .A(\u_div/PartRem[2][5] ), .B(\u_div/u_add_PartRem_2_1/n2 ), .Y(
        \u_div/CryTmp[1][6] ) );
  OR2X2 U42 ( .A(\u_div/PartRem[9][5] ), .B(\u_div/u_add_PartRem_2_8/n2 ), .Y(
        \u_div/CryTmp[8][6] ) );
  OR2X2 U43 ( .A(\u_div/PartRem[37][5] ), .B(\u_div/u_add_PartRem_2_36/n2 ), 
        .Y(\u_div/CryTmp[36][6] ) );
  NOR2BX2 U44 ( .AN(\u_div/PartRem[64][0] ), .B(n8), .Y(\u_div/CryTmp[59][6] )
         );
  MXI2X1 U45 ( .A(\u_div/SumTmp[1][1] ), .B(\u_div/SumTmp[1][1] ), .S0(
        \u_div/CryTmp[1][6] ), .Y(n1) );
  OR2X2 U46 ( .A(\u_div/PartRem[47][5] ), .B(\u_div/u_add_PartRem_2_46/n2 ), 
        .Y(\u_div/CryTmp[46][6] ) );
  ADDHX2 U47 ( .A(\u_div/PartRem[37][4] ), .B(\u_div/u_add_PartRem_2_36/n3 ), 
        .CO(\u_div/u_add_PartRem_2_36/n2 ), .S(\u_div/SumTmp[36][4] ) );
  OR2X8 U48 ( .A(\u_div/PartRem[27][5] ), .B(\u_div/u_add_PartRem_2_26/n2 ), 
        .Y(\u_div/CryTmp[26][6] ) );
  ADDHX2 U49 ( .A(\u_div/PartRem[27][4] ), .B(\u_div/u_add_PartRem_2_26/n3 ), 
        .CO(\u_div/u_add_PartRem_2_26/n2 ), .S(\u_div/SumTmp[26][4] ) );
  ADDHX2 U50 ( .A(\u_div/PartRem[19][4] ), .B(\u_div/u_add_PartRem_2_18/n3 ), 
        .CO(\u_div/u_add_PartRem_2_18/n2 ), .S(\u_div/SumTmp[18][4] ) );
  XOR2XL U51 ( .A(\u_div/CryTmp[8][6] ), .B(n3), .Y(\u_div/QInv[8] ) );
  MXI2X4 U52 ( .A(\u_div/SumTmp[8][2] ), .B(\u_div/PartRem[9][2] ), .S0(
        \u_div/CryTmp[8][6] ), .Y(\u_div/PartRem[8][3] ) );
  OR2X6 U53 ( .A(\u_div/PartRem[59][2] ), .B(\u_div/PartRem[59][3] ), .Y(
        \u_div/u_add_PartRem_2_58/n3 ) );
  XOR2X1 U54 ( .A(\u_div/CryTmp[0][6] ), .B(n5), .Y(\u_div/QInv[0] ) );
  AO21X1 U55 ( .A0(\u_div/PartRem[1][4] ), .A1(n6), .B0(\u_div/PartRem[1][5] ), 
        .Y(\u_div/CryTmp[0][6] ) );
  ADDHXL U56 ( .A(\u_div/PartRem[58][4] ), .B(\u_div/u_add_PartRem_2_57/n3 ), 
        .CO(\u_div/u_add_PartRem_2_57/n2 ), .S(\u_div/SumTmp[57][4] ) );
  ADDHXL U57 ( .A(\u_div/PartRem[57][4] ), .B(\u_div/u_add_PartRem_2_56/n3 ), 
        .CO(\u_div/u_add_PartRem_2_56/n2 ), .S(\u_div/SumTmp[56][4] ) );
  ADDHXL U58 ( .A(\u_div/PartRem[56][4] ), .B(\u_div/u_add_PartRem_2_55/n3 ), 
        .CO(\u_div/u_add_PartRem_2_55/n2 ), .S(\u_div/SumTmp[55][4] ) );
  ADDHXL U59 ( .A(\u_div/PartRem[54][4] ), .B(\u_div/u_add_PartRem_2_53/n3 ), 
        .CO(\u_div/u_add_PartRem_2_53/n2 ), .S(\u_div/SumTmp[53][4] ) );
  ADDHXL U60 ( .A(\u_div/PartRem[49][4] ), .B(\u_div/u_add_PartRem_2_48/n3 ), 
        .CO(\u_div/u_add_PartRem_2_48/n2 ), .S(\u_div/SumTmp[48][4] ) );
  ADDHXL U61 ( .A(\u_div/PartRem[47][4] ), .B(\u_div/u_add_PartRem_2_46/n3 ), 
        .CO(\u_div/u_add_PartRem_2_46/n2 ), .S(\u_div/SumTmp[46][4] ) );
  ADDHXL U62 ( .A(\u_div/PartRem[45][4] ), .B(\u_div/u_add_PartRem_2_44/n3 ), 
        .CO(\u_div/u_add_PartRem_2_44/n2 ), .S(\u_div/SumTmp[44][4] ) );
  ADDHXL U63 ( .A(\u_div/PartRem[39][4] ), .B(\u_div/u_add_PartRem_2_38/n3 ), 
        .CO(\u_div/u_add_PartRem_2_38/n2 ), .S(\u_div/SumTmp[38][4] ) );
  ADDHXL U64 ( .A(\u_div/PartRem[35][4] ), .B(\u_div/u_add_PartRem_2_34/n3 ), 
        .CO(\u_div/u_add_PartRem_2_34/n2 ), .S(\u_div/SumTmp[34][4] ) );
  ADDHXL U65 ( .A(\u_div/PartRem[34][4] ), .B(\u_div/u_add_PartRem_2_33/n3 ), 
        .CO(\u_div/u_add_PartRem_2_33/n2 ), .S(\u_div/SumTmp[33][4] ) );
  ADDHXL U66 ( .A(\u_div/PartRem[32][4] ), .B(\u_div/u_add_PartRem_2_31/n3 ), 
        .CO(\u_div/u_add_PartRem_2_31/n2 ), .S(\u_div/SumTmp[31][4] ) );
  ADDHXL U67 ( .A(\u_div/PartRem[29][4] ), .B(\u_div/u_add_PartRem_2_28/n3 ), 
        .CO(\u_div/u_add_PartRem_2_28/n2 ), .S(\u_div/SumTmp[28][4] ) );
  ADDHXL U68 ( .A(\u_div/PartRem[25][4] ), .B(\u_div/u_add_PartRem_2_24/n3 ), 
        .CO(\u_div/u_add_PartRem_2_24/n2 ), .S(\u_div/SumTmp[24][4] ) );
  ADDHXL U69 ( .A(\u_div/PartRem[24][4] ), .B(\u_div/u_add_PartRem_2_23/n3 ), 
        .CO(\u_div/u_add_PartRem_2_23/n2 ), .S(\u_div/SumTmp[23][4] ) );
  ADDHXL U70 ( .A(\u_div/PartRem[22][4] ), .B(\u_div/u_add_PartRem_2_21/n3 ), 
        .CO(\u_div/u_add_PartRem_2_21/n2 ), .S(\u_div/SumTmp[21][4] ) );
  ADDHXL U71 ( .A(\u_div/PartRem[17][4] ), .B(\u_div/u_add_PartRem_2_16/n3 ), 
        .CO(\u_div/u_add_PartRem_2_16/n2 ), .S(\u_div/SumTmp[16][4] ) );
  ADDHXL U72 ( .A(\u_div/PartRem[15][4] ), .B(\u_div/u_add_PartRem_2_14/n3 ), 
        .CO(\u_div/u_add_PartRem_2_14/n2 ), .S(\u_div/SumTmp[14][4] ) );
  ADDHXL U73 ( .A(\u_div/PartRem[9][4] ), .B(\u_div/u_add_PartRem_2_8/n3 ), 
        .CO(\u_div/u_add_PartRem_2_8/n2 ), .S(\u_div/SumTmp[8][4] ) );
  ADDHXL U74 ( .A(\u_div/PartRem[7][4] ), .B(\u_div/u_add_PartRem_2_6/n3 ), 
        .CO(\u_div/u_add_PartRem_2_6/n2 ), .S(\u_div/SumTmp[6][4] ) );
  ADDHXL U75 ( .A(\u_div/PartRem[2][4] ), .B(\u_div/u_add_PartRem_2_1/n3 ), 
        .CO(\u_div/u_add_PartRem_2_1/n2 ), .S(\u_div/SumTmp[1][4] ) );
  ADDHXL U76 ( .A(\u_div/PartRem[55][4] ), .B(\u_div/u_add_PartRem_2_54/n3 ), 
        .CO(\u_div/u_add_PartRem_2_54/n2 ), .S(\u_div/SumTmp[54][4] ) );
  ADDHXL U77 ( .A(\u_div/PartRem[50][4] ), .B(\u_div/u_add_PartRem_2_49/n3 ), 
        .CO(\u_div/u_add_PartRem_2_49/n2 ), .S(\u_div/SumTmp[49][4] ) );
  ADDHXL U78 ( .A(\u_div/PartRem[44][4] ), .B(\u_div/u_add_PartRem_2_43/n3 ), 
        .CO(\u_div/u_add_PartRem_2_43/n2 ), .S(\u_div/SumTmp[43][4] ) );
  ADDHXL U79 ( .A(\u_div/PartRem[42][4] ), .B(\u_div/u_add_PartRem_2_41/n3 ), 
        .CO(\u_div/u_add_PartRem_2_41/n2 ), .S(\u_div/SumTmp[41][4] ) );
  ADDHXL U80 ( .A(\u_div/PartRem[40][4] ), .B(\u_div/u_add_PartRem_2_39/n3 ), 
        .CO(\u_div/u_add_PartRem_2_39/n2 ), .S(\u_div/SumTmp[39][4] ) );
  ADDHXL U81 ( .A(\u_div/PartRem[30][4] ), .B(\u_div/u_add_PartRem_2_29/n3 ), 
        .CO(\u_div/u_add_PartRem_2_29/n2 ), .S(\u_div/SumTmp[29][4] ) );
  ADDHXL U82 ( .A(\u_div/PartRem[21][4] ), .B(\u_div/u_add_PartRem_2_20/n3 ), 
        .CO(\u_div/u_add_PartRem_2_20/n2 ), .S(\u_div/SumTmp[20][4] ) );
  ADDHXL U83 ( .A(\u_div/PartRem[16][4] ), .B(\u_div/u_add_PartRem_2_15/n3 ), 
        .CO(\u_div/u_add_PartRem_2_15/n2 ), .S(\u_div/SumTmp[15][4] ) );
  ADDHXL U84 ( .A(\u_div/PartRem[12][4] ), .B(\u_div/u_add_PartRem_2_11/n3 ), 
        .CO(\u_div/u_add_PartRem_2_11/n2 ), .S(\u_div/SumTmp[11][4] ) );
  ADDHXL U85 ( .A(\u_div/PartRem[11][4] ), .B(\u_div/u_add_PartRem_2_10/n3 ), 
        .CO(\u_div/u_add_PartRem_2_10/n2 ), .S(\u_div/SumTmp[10][4] ) );
  ADDHXL U86 ( .A(\u_div/PartRem[10][4] ), .B(\u_div/u_add_PartRem_2_9/n3 ), 
        .CO(\u_div/u_add_PartRem_2_9/n2 ), .S(\u_div/SumTmp[9][4] ) );
  ADDHXL U87 ( .A(\u_div/PartRem[6][4] ), .B(\u_div/u_add_PartRem_2_5/n3 ), 
        .CO(\u_div/u_add_PartRem_2_5/n2 ), .S(\u_div/SumTmp[5][4] ) );
  ADDHXL U88 ( .A(\u_div/PartRem[20][4] ), .B(\u_div/u_add_PartRem_2_19/n3 ), 
        .CO(\u_div/u_add_PartRem_2_19/n2 ), .S(\u_div/SumTmp[19][4] ) );
  ADDHXL U89 ( .A(\u_div/PartRem[36][4] ), .B(\u_div/u_add_PartRem_2_35/n3 ), 
        .CO(\u_div/u_add_PartRem_2_35/n2 ), .S(\u_div/SumTmp[35][4] ) );
  ADDHXL U90 ( .A(\u_div/PartRem[26][4] ), .B(\u_div/u_add_PartRem_2_25/n3 ), 
        .CO(\u_div/u_add_PartRem_2_25/n2 ), .S(\u_div/SumTmp[25][4] ) );
  ADDHXL U91 ( .A(\u_div/PartRem[31][4] ), .B(\u_div/u_add_PartRem_2_30/n3 ), 
        .CO(\u_div/u_add_PartRem_2_30/n2 ), .S(\u_div/SumTmp[30][4] ) );
  ADDHXL U92 ( .A(\u_div/PartRem[41][4] ), .B(\u_div/u_add_PartRem_2_40/n3 ), 
        .CO(\u_div/u_add_PartRem_2_40/n2 ), .S(\u_div/SumTmp[40][4] ) );
  ADDHXL U93 ( .A(\u_div/PartRem[46][4] ), .B(\u_div/u_add_PartRem_2_45/n3 ), 
        .CO(\u_div/u_add_PartRem_2_45/n2 ), .S(\u_div/SumTmp[45][4] ) );
  ADDHXL U94 ( .A(\u_div/PartRem[51][4] ), .B(\u_div/u_add_PartRem_2_50/n3 ), 
        .CO(\u_div/u_add_PartRem_2_50/n2 ), .S(\u_div/SumTmp[50][4] ) );
  MXI2X2 U95 ( .A(\u_div/SumTmp[18][2] ), .B(\u_div/PartRem[19][2] ), .S0(
        \u_div/CryTmp[18][6] ), .Y(\u_div/PartRem[18][3] ) );
  MXI2X2 U96 ( .A(\u_div/SumTmp[26][2] ), .B(\u_div/PartRem[27][2] ), .S0(
        \u_div/CryTmp[26][6] ), .Y(\u_div/PartRem[26][3] ) );
  MXI2X2 U97 ( .A(\u_div/SumTmp[36][2] ), .B(\u_div/PartRem[37][2] ), .S0(
        \u_div/CryTmp[36][6] ), .Y(\u_div/PartRem[36][3] ) );
  MXI2X2 U98 ( .A(\u_div/SumTmp[46][2] ), .B(\u_div/PartRem[47][2] ), .S0(
        \u_div/CryTmp[46][6] ), .Y(\u_div/PartRem[46][3] ) );
  MXI2X2 U99 ( .A(\u_div/SumTmp[13][2] ), .B(\u_div/PartRem[14][2] ), .S0(
        \u_div/CryTmp[13][6] ), .Y(\u_div/PartRem[13][3] ) );
  MXI2X2 U100 ( .A(\u_div/SumTmp[51][2] ), .B(\u_div/PartRem[52][2] ), .S0(
        \u_div/CryTmp[51][6] ), .Y(\u_div/PartRem[51][3] ) );
  MXI2X2 U101 ( .A(\u_div/SumTmp[4][2] ), .B(\u_div/PartRem[5][2] ), .S0(
        \u_div/CryTmp[4][6] ), .Y(\u_div/PartRem[4][3] ) );
  OR2X2 U102 ( .A(\u_div/PartRem[24][2] ), .B(\u_div/PartRem[24][3] ), .Y(
        \u_div/u_add_PartRem_2_23/n3 ) );
  OR2X2 U103 ( .A(\u_div/PartRem[22][2] ), .B(\u_div/PartRem[22][3] ), .Y(
        \u_div/u_add_PartRem_2_21/n3 ) );
  OR2X2 U104 ( .A(\u_div/PartRem[21][2] ), .B(\u_div/PartRem[21][3] ), .Y(
        \u_div/u_add_PartRem_2_20/n3 ) );
  OR2X2 U105 ( .A(\u_div/PartRem[14][2] ), .B(\u_div/PartRem[14][3] ), .Y(
        \u_div/u_add_PartRem_2_13/n3 ) );
  OR2X2 U106 ( .A(\u_div/PartRem[10][2] ), .B(\u_div/PartRem[10][3] ), .Y(
        \u_div/u_add_PartRem_2_9/n3 ) );
  OR2X2 U107 ( .A(\u_div/PartRem[20][2] ), .B(\u_div/PartRem[20][3] ), .Y(
        \u_div/u_add_PartRem_2_19/n3 ) );
  OR2X2 U108 ( .A(\u_div/PartRem[19][2] ), .B(\u_div/PartRem[19][3] ), .Y(
        \u_div/u_add_PartRem_2_18/n3 ) );
  OR2X2 U109 ( .A(\u_div/PartRem[27][2] ), .B(\u_div/PartRem[27][3] ), .Y(
        \u_div/u_add_PartRem_2_26/n3 ) );
  OR2X2 U110 ( .A(\u_div/PartRem[9][2] ), .B(\u_div/PartRem[9][3] ), .Y(
        \u_div/u_add_PartRem_2_8/n3 ) );
  OR2X2 U111 ( .A(\u_div/PartRem[30][2] ), .B(\u_div/PartRem[30][3] ), .Y(
        \u_div/u_add_PartRem_2_29/n3 ) );
  OR2X2 U112 ( .A(\u_div/PartRem[37][2] ), .B(\u_div/PartRem[37][3] ), .Y(
        \u_div/u_add_PartRem_2_36/n3 ) );
  OR2X2 U113 ( .A(\u_div/PartRem[40][2] ), .B(\u_div/PartRem[40][3] ), .Y(
        \u_div/u_add_PartRem_2_39/n3 ) );
  OR2X2 U114 ( .A(\u_div/PartRem[47][2] ), .B(\u_div/PartRem[47][3] ), .Y(
        \u_div/u_add_PartRem_2_46/n3 ) );
  OR2X2 U115 ( .A(\u_div/PartRem[2][2] ), .B(\u_div/PartRem[2][3] ), .Y(
        \u_div/u_add_PartRem_2_1/n3 ) );
  OR2X2 U116 ( .A(\u_div/PartRem[56][2] ), .B(\u_div/PartRem[56][3] ), .Y(
        \u_div/u_add_PartRem_2_55/n3 ) );
  ADDHX2 U117 ( .A(\u_div/PartRem[59][4] ), .B(\u_div/u_add_PartRem_2_58/n3 ), 
        .CO(\u_div/u_add_PartRem_2_58/n2 ), .S(\u_div/SumTmp[58][4] ) );
  ADDHX1 U118 ( .A(\u_div/PartRem[4][4] ), .B(\u_div/u_add_PartRem_2_3/n3 ), 
        .CO(\u_div/u_add_PartRem_2_3/n2 ), .S(\u_div/SumTmp[3][4] ) );
  NAND2BX2 U119 ( .AN(\u_div/PartRem[1][3] ), .B(n1), .Y(n6) );
  OR2X1 U120 ( .A(\u_div/PartRem[53][2] ), .B(\u_div/PartRem[53][3] ), .Y(
        \u_div/u_add_PartRem_2_52/n3 ) );
  OR2X1 U121 ( .A(\u_div/PartRem[48][2] ), .B(\u_div/PartRem[48][3] ), .Y(
        \u_div/u_add_PartRem_2_47/n3 ) );
  OR2X1 U122 ( .A(\u_div/PartRem[43][2] ), .B(\u_div/PartRem[43][3] ), .Y(
        \u_div/u_add_PartRem_2_42/n3 ) );
  OR2X1 U123 ( .A(\u_div/PartRem[38][2] ), .B(\u_div/PartRem[38][3] ), .Y(
        \u_div/u_add_PartRem_2_37/n3 ) );
  OR2X1 U124 ( .A(\u_div/PartRem[33][2] ), .B(\u_div/PartRem[33][3] ), .Y(
        \u_div/u_add_PartRem_2_32/n3 ) );
  OR2X1 U125 ( .A(\u_div/PartRem[28][2] ), .B(\u_div/PartRem[28][3] ), .Y(
        \u_div/u_add_PartRem_2_27/n3 ) );
  OR2X1 U126 ( .A(\u_div/PartRem[23][2] ), .B(\u_div/PartRem[23][3] ), .Y(
        \u_div/u_add_PartRem_2_22/n3 ) );
  XNOR2XL U127 ( .A(\u_div/PartRem[64][0] ), .B(n8), .Y(\u_div/SumTmp[59][4] )
         );
  XOR2XL U128 ( .A(\u_div/CryTmp[55][6] ), .B(n5), .Y(\u_div/QInv[55] ) );
  XOR2XL U129 ( .A(\u_div/CryTmp[44][6] ), .B(n5), .Y(\u_div/QInv[44] ) );
  XOR2XL U130 ( .A(\u_div/CryTmp[41][6] ), .B(n5), .Y(\u_div/QInv[41] ) );
  XOR2XL U131 ( .A(\u_div/CryTmp[31][6] ), .B(n5), .Y(\u_div/QInv[31] ) );
  XOR2XL U132 ( .A(\u_div/CryTmp[20][6] ), .B(n5), .Y(\u_div/QInv[20] ) );
  XOR2XL U133 ( .A(\u_div/CryTmp[12][6] ), .B(n5), .Y(\u_div/QInv[12] ) );
  XOR2XL U134 ( .A(\u_div/CryTmp[11][6] ), .B(n4), .Y(\u_div/QInv[11] ) );
  XOR2XL U135 ( .A(\u_div/CryTmp[50][6] ), .B(n3), .Y(\u_div/QInv[50] ) );
  XOR2XL U136 ( .A(\u_div/CryTmp[51][6] ), .B(n4), .Y(\u_div/QInv[51] ) );
  XOR2XL U137 ( .A(\u_div/CryTmp[43][6] ), .B(n4), .Y(\u_div/QInv[43] ) );
  XOR2XL U138 ( .A(\u_div/CryTmp[42][6] ), .B(n3), .Y(\u_div/QInv[42] ) );
  XOR2XL U139 ( .A(\u_div/CryTmp[40][6] ), .B(n4), .Y(\u_div/QInv[40] ) );
  XOR2XL U140 ( .A(\u_div/CryTmp[30][6] ), .B(n4), .Y(\u_div/QInv[30] ) );
  XOR2XL U141 ( .A(\u_div/CryTmp[21][6] ), .B(n3), .Y(\u_div/QInv[21] ) );
  XOR2XL U142 ( .A(\u_div/CryTmp[16][6] ), .B(n5), .Y(\u_div/QInv[16] ) );
  XOR2XL U143 ( .A(\u_div/CryTmp[13][6] ), .B(n4), .Y(\u_div/QInv[13] ) );
  XOR2XL U144 ( .A(\u_div/CryTmp[4][6] ), .B(n5), .Y(\u_div/QInv[4] ) );
  XOR2XL U145 ( .A(\u_div/CryTmp[5][6] ), .B(n4), .Y(\u_div/QInv[5] ) );
  XOR2XL U146 ( .A(\u_div/CryTmp[6][6] ), .B(n5), .Y(\u_div/QInv[6] ) );
  XOR2XL U147 ( .A(\u_div/CryTmp[10][6] ), .B(n5), .Y(\u_div/QInv[10] ) );
  XOR2XL U148 ( .A(\u_div/CryTmp[3][6] ), .B(n3), .Y(\u_div/QInv[3] ) );
  INVXL U149 ( .A(\u_div/PartRem[59][2] ), .Y(\u_div/SumTmp[58][2] ) );
  INVXL U150 ( .A(\u_div/PartRem[53][2] ), .Y(\u_div/SumTmp[52][2] ) );
  INVXL U151 ( .A(\u_div/PartRem[48][2] ), .Y(\u_div/SumTmp[47][2] ) );
  INVXL U152 ( .A(\u_div/PartRem[43][2] ), .Y(\u_div/SumTmp[42][2] ) );
  INVXL U153 ( .A(\u_div/PartRem[38][2] ), .Y(\u_div/SumTmp[37][2] ) );
  INVXL U154 ( .A(\u_div/PartRem[33][2] ), .Y(\u_div/SumTmp[32][2] ) );
  INVXL U155 ( .A(\u_div/PartRem[28][2] ), .Y(\u_div/SumTmp[27][2] ) );
  INVXL U156 ( .A(\u_div/PartRem[23][2] ), .Y(\u_div/SumTmp[22][2] ) );
  INVXL U157 ( .A(\u_div/PartRem[20][2] ), .Y(\u_div/SumTmp[19][2] ) );
  INVX3 U158 ( .A(n2), .Y(n3) );
  CLKINVX1 U159 ( .A(\u_div/QInv[63] ), .Y(n2) );
  OR2X1 U160 ( .A(\u_div/PartRem[18][2] ), .B(\u_div/PartRem[18][3] ), .Y(
        \u_div/u_add_PartRem_2_17/n3 ) );
  OR2X1 U161 ( .A(\u_div/PartRem[13][2] ), .B(\u_div/PartRem[13][3] ), .Y(
        \u_div/u_add_PartRem_2_12/n3 ) );
  OR2X1 U162 ( .A(\u_div/PartRem[8][2] ), .B(\u_div/PartRem[8][3] ), .Y(
        \u_div/u_add_PartRem_2_7/n3 ) );
  OR2X1 U163 ( .A(\u_div/PartRem[3][2] ), .B(\u_div/PartRem[3][3] ), .Y(
        \u_div/u_add_PartRem_2_2/n3 ) );
  MXI2X1 U164 ( .A(\u_div/SumTmp[56][2] ), .B(\u_div/PartRem[57][2] ), .S0(
        \u_div/CryTmp[56][6] ), .Y(\u_div/PartRem[56][3] ) );
  CLKINVX1 U165 ( .A(\u_div/PartRem[57][2] ), .Y(\u_div/SumTmp[56][2] ) );
  MXI2X1 U166 ( .A(\u_div/SumTmp[19][2] ), .B(\u_div/PartRem[20][2] ), .S0(
        \u_div/CryTmp[19][6] ), .Y(\u_div/PartRem[19][3] ) );
  MXI2X1 U167 ( .A(\u_div/SumTmp[16][2] ), .B(\u_div/PartRem[17][2] ), .S0(
        \u_div/CryTmp[16][6] ), .Y(\u_div/PartRem[16][3] ) );
  CLKINVX1 U168 ( .A(\u_div/PartRem[17][2] ), .Y(\u_div/SumTmp[16][2] ) );
  MXI2X1 U169 ( .A(\u_div/SumTmp[12][2] ), .B(\u_div/PartRem[13][2] ), .S0(
        \u_div/CryTmp[12][6] ), .Y(\u_div/PartRem[12][3] ) );
  CLKINVX1 U170 ( .A(\u_div/PartRem[13][2] ), .Y(\u_div/SumTmp[12][2] ) );
  MXI2X1 U171 ( .A(\u_div/SumTmp[9][2] ), .B(\u_div/PartRem[10][2] ), .S0(
        \u_div/CryTmp[9][6] ), .Y(\u_div/PartRem[9][3] ) );
  CLKINVX1 U172 ( .A(\u_div/PartRem[10][2] ), .Y(\u_div/SumTmp[9][2] ) );
  MXI2X1 U173 ( .A(\u_div/SumTmp[6][2] ), .B(\u_div/PartRem[7][2] ), .S0(
        \u_div/CryTmp[6][6] ), .Y(\u_div/PartRem[6][3] ) );
  CLKINVX1 U174 ( .A(\u_div/PartRem[7][2] ), .Y(\u_div/SumTmp[6][2] ) );
  CLKINVX1 U175 ( .A(\u_div/PartRem[3][2] ), .Y(\u_div/SumTmp[2][2] ) );
  MXI2X1 U176 ( .A(n7), .B(\u_div/PartRem[62][0] ), .S0(\u_div/CryTmp[59][6] ), 
        .Y(\u_div/PartRem[59][3] ) );
  CLKINVX1 U177 ( .A(\u_div/PartRem[62][0] ), .Y(n7) );
  CLKINVX1 U178 ( .A(\u_div/PartRem[4][2] ), .Y(\u_div/SumTmp[3][2] ) );
  CLKINVX1 U179 ( .A(\u_div/PartRem[19][2] ), .Y(\u_div/SumTmp[18][2] ) );
  CLKINVX1 U180 ( .A(\u_div/PartRem[14][2] ), .Y(\u_div/SumTmp[13][2] ) );
  CLKINVX1 U181 ( .A(\u_div/PartRem[9][2] ), .Y(\u_div/SumTmp[8][2] ) );
  MXI2X1 U182 ( .A(\u_div/SumTmp[58][2] ), .B(\u_div/PartRem[59][2] ), .S0(
        \u_div/CryTmp[58][6] ), .Y(\u_div/PartRem[58][3] ) );
  MXI2X1 U183 ( .A(\u_div/SumTmp[57][2] ), .B(\u_div/PartRem[58][2] ), .S0(
        \u_div/CryTmp[57][6] ), .Y(\u_div/PartRem[57][3] ) );
  CLKINVX1 U184 ( .A(\u_div/PartRem[58][2] ), .Y(\u_div/SumTmp[57][2] ) );
  MXI2X1 U185 ( .A(\u_div/SumTmp[54][2] ), .B(\u_div/PartRem[55][2] ), .S0(
        \u_div/CryTmp[54][6] ), .Y(\u_div/PartRem[54][3] ) );
  CLKINVX1 U186 ( .A(\u_div/PartRem[55][2] ), .Y(\u_div/SumTmp[54][2] ) );
  MXI2X1 U187 ( .A(\u_div/SumTmp[55][2] ), .B(\u_div/PartRem[56][2] ), .S0(
        \u_div/CryTmp[55][6] ), .Y(\u_div/PartRem[55][3] ) );
  CLKINVX1 U188 ( .A(\u_div/PartRem[56][2] ), .Y(\u_div/SumTmp[55][2] ) );
  MXI2X1 U189 ( .A(\u_div/SumTmp[52][2] ), .B(\u_div/PartRem[53][2] ), .S0(
        \u_div/CryTmp[52][6] ), .Y(\u_div/PartRem[52][3] ) );
  CLKINVX1 U190 ( .A(\u_div/PartRem[52][2] ), .Y(\u_div/SumTmp[51][2] ) );
  MXI2X1 U191 ( .A(\u_div/SumTmp[49][2] ), .B(\u_div/PartRem[50][2] ), .S0(
        \u_div/CryTmp[49][6] ), .Y(\u_div/PartRem[49][3] ) );
  CLKINVX1 U192 ( .A(\u_div/PartRem[50][2] ), .Y(\u_div/SumTmp[49][2] ) );
  MXI2X1 U193 ( .A(\u_div/SumTmp[50][2] ), .B(\u_div/PartRem[51][2] ), .S0(
        \u_div/CryTmp[50][6] ), .Y(\u_div/PartRem[50][3] ) );
  CLKINVX1 U194 ( .A(\u_div/PartRem[51][2] ), .Y(\u_div/SumTmp[50][2] ) );
  MXI2X1 U195 ( .A(\u_div/SumTmp[47][2] ), .B(\u_div/PartRem[48][2] ), .S0(
        \u_div/CryTmp[47][6] ), .Y(\u_div/PartRem[47][3] ) );
  CLKINVX1 U196 ( .A(\u_div/PartRem[47][2] ), .Y(\u_div/SumTmp[46][2] ) );
  MXI2X1 U197 ( .A(\u_div/SumTmp[44][2] ), .B(\u_div/PartRem[45][2] ), .S0(
        \u_div/CryTmp[44][6] ), .Y(\u_div/PartRem[44][3] ) );
  CLKINVX1 U198 ( .A(\u_div/PartRem[45][2] ), .Y(\u_div/SumTmp[44][2] ) );
  MXI2X1 U199 ( .A(\u_div/SumTmp[45][2] ), .B(\u_div/PartRem[46][2] ), .S0(
        \u_div/CryTmp[45][6] ), .Y(\u_div/PartRem[45][3] ) );
  CLKINVX1 U200 ( .A(\u_div/PartRem[46][2] ), .Y(\u_div/SumTmp[45][2] ) );
  MXI2X1 U201 ( .A(\u_div/SumTmp[42][2] ), .B(\u_div/PartRem[43][2] ), .S0(
        \u_div/CryTmp[42][6] ), .Y(\u_div/PartRem[42][3] ) );
  CLKINVX1 U202 ( .A(\u_div/PartRem[42][2] ), .Y(\u_div/SumTmp[41][2] ) );
  MXI2X1 U203 ( .A(\u_div/SumTmp[39][2] ), .B(\u_div/PartRem[40][2] ), .S0(
        \u_div/CryTmp[39][6] ), .Y(\u_div/PartRem[39][3] ) );
  CLKINVX1 U204 ( .A(\u_div/PartRem[40][2] ), .Y(\u_div/SumTmp[39][2] ) );
  MXI2X1 U205 ( .A(\u_div/SumTmp[40][2] ), .B(\u_div/PartRem[41][2] ), .S0(
        \u_div/CryTmp[40][6] ), .Y(\u_div/PartRem[40][3] ) );
  CLKINVX1 U206 ( .A(\u_div/PartRem[41][2] ), .Y(\u_div/SumTmp[40][2] ) );
  MXI2X1 U207 ( .A(\u_div/SumTmp[37][2] ), .B(\u_div/PartRem[38][2] ), .S0(
        \u_div/CryTmp[37][6] ), .Y(\u_div/PartRem[37][3] ) );
  CLKINVX1 U208 ( .A(\u_div/PartRem[37][2] ), .Y(\u_div/SumTmp[36][2] ) );
  MXI2X1 U209 ( .A(\u_div/SumTmp[34][2] ), .B(\u_div/PartRem[35][2] ), .S0(
        \u_div/CryTmp[34][6] ), .Y(\u_div/PartRem[34][3] ) );
  CLKINVX1 U210 ( .A(\u_div/PartRem[35][2] ), .Y(\u_div/SumTmp[34][2] ) );
  MXI2X1 U211 ( .A(\u_div/SumTmp[35][2] ), .B(\u_div/PartRem[36][2] ), .S0(
        \u_div/CryTmp[35][6] ), .Y(\u_div/PartRem[35][3] ) );
  CLKINVX1 U212 ( .A(\u_div/PartRem[36][2] ), .Y(\u_div/SumTmp[35][2] ) );
  MXI2X1 U213 ( .A(\u_div/SumTmp[32][2] ), .B(\u_div/PartRem[33][2] ), .S0(
        \u_div/CryTmp[32][6] ), .Y(\u_div/PartRem[32][3] ) );
  CLKINVX1 U214 ( .A(\u_div/PartRem[32][2] ), .Y(\u_div/SumTmp[31][2] ) );
  MXI2X1 U215 ( .A(\u_div/SumTmp[29][2] ), .B(\u_div/PartRem[30][2] ), .S0(
        \u_div/CryTmp[29][6] ), .Y(\u_div/PartRem[29][3] ) );
  CLKINVX1 U216 ( .A(\u_div/PartRem[30][2] ), .Y(\u_div/SumTmp[29][2] ) );
  MXI2X1 U217 ( .A(\u_div/SumTmp[30][2] ), .B(\u_div/PartRem[31][2] ), .S0(
        \u_div/CryTmp[30][6] ), .Y(\u_div/PartRem[30][3] ) );
  CLKINVX1 U218 ( .A(\u_div/PartRem[31][2] ), .Y(\u_div/SumTmp[30][2] ) );
  MXI2X1 U219 ( .A(\u_div/SumTmp[27][2] ), .B(\u_div/PartRem[28][2] ), .S0(
        \u_div/CryTmp[27][6] ), .Y(\u_div/PartRem[27][3] ) );
  CLKINVX1 U220 ( .A(\u_div/PartRem[27][2] ), .Y(\u_div/SumTmp[26][2] ) );
  MXI2X1 U221 ( .A(\u_div/SumTmp[24][2] ), .B(\u_div/PartRem[25][2] ), .S0(
        \u_div/CryTmp[24][6] ), .Y(\u_div/PartRem[24][3] ) );
  CLKINVX1 U222 ( .A(\u_div/PartRem[25][2] ), .Y(\u_div/SumTmp[24][2] ) );
  MXI2X1 U223 ( .A(\u_div/SumTmp[25][2] ), .B(\u_div/PartRem[26][2] ), .S0(
        \u_div/CryTmp[25][6] ), .Y(\u_div/PartRem[25][3] ) );
  CLKINVX1 U224 ( .A(\u_div/PartRem[26][2] ), .Y(\u_div/SumTmp[25][2] ) );
  MXI2X1 U225 ( .A(\u_div/SumTmp[22][2] ), .B(\u_div/PartRem[23][2] ), .S0(
        \u_div/CryTmp[22][6] ), .Y(\u_div/PartRem[22][3] ) );
  MXI2X1 U226 ( .A(\u_div/SumTmp[21][2] ), .B(\u_div/PartRem[22][2] ), .S0(
        \u_div/CryTmp[21][6] ), .Y(\u_div/PartRem[21][3] ) );
  CLKINVX1 U227 ( .A(\u_div/PartRem[22][2] ), .Y(\u_div/SumTmp[21][2] ) );
  MXI2X1 U228 ( .A(\u_div/SumTmp[17][2] ), .B(\u_div/PartRem[18][2] ), .S0(
        \u_div/CryTmp[17][6] ), .Y(\u_div/PartRem[17][3] ) );
  CLKINVX1 U229 ( .A(\u_div/PartRem[18][2] ), .Y(\u_div/SumTmp[17][2] ) );
  MXI2X1 U230 ( .A(\u_div/SumTmp[15][2] ), .B(\u_div/PartRem[16][2] ), .S0(
        \u_div/CryTmp[15][6] ), .Y(\u_div/PartRem[15][3] ) );
  CLKINVX1 U231 ( .A(\u_div/PartRem[16][2] ), .Y(\u_div/SumTmp[15][2] ) );
  MXI2X1 U232 ( .A(\u_div/SumTmp[14][2] ), .B(\u_div/PartRem[15][2] ), .S0(
        \u_div/CryTmp[14][6] ), .Y(\u_div/PartRem[14][3] ) );
  CLKINVX1 U233 ( .A(\u_div/PartRem[15][2] ), .Y(\u_div/SumTmp[14][2] ) );
  MXI2X1 U234 ( .A(\u_div/SumTmp[11][2] ), .B(\u_div/PartRem[12][2] ), .S0(
        \u_div/CryTmp[11][6] ), .Y(\u_div/PartRem[11][3] ) );
  CLKINVX1 U235 ( .A(\u_div/PartRem[12][2] ), .Y(\u_div/SumTmp[11][2] ) );
  MXI2X1 U236 ( .A(\u_div/SumTmp[10][2] ), .B(\u_div/PartRem[11][2] ), .S0(
        \u_div/CryTmp[10][6] ), .Y(\u_div/PartRem[10][3] ) );
  CLKINVX1 U237 ( .A(\u_div/PartRem[11][2] ), .Y(\u_div/SumTmp[10][2] ) );
  MXI2X1 U238 ( .A(\u_div/SumTmp[7][2] ), .B(\u_div/PartRem[8][2] ), .S0(
        \u_div/CryTmp[7][6] ), .Y(\u_div/PartRem[7][3] ) );
  CLKINVX1 U239 ( .A(\u_div/PartRem[8][2] ), .Y(\u_div/SumTmp[7][2] ) );
  MXI2X1 U240 ( .A(\u_div/SumTmp[5][2] ), .B(\u_div/PartRem[6][2] ), .S0(
        \u_div/CryTmp[5][6] ), .Y(\u_div/PartRem[5][3] ) );
  CLKINVX1 U241 ( .A(\u_div/PartRem[6][2] ), .Y(\u_div/SumTmp[5][2] ) );
  CLKINVX1 U242 ( .A(\u_div/PartRem[5][2] ), .Y(\u_div/SumTmp[4][2] ) );
  MXI2X1 U243 ( .A(\u_div/SumTmp[53][2] ), .B(\u_div/PartRem[54][2] ), .S0(
        \u_div/CryTmp[53][6] ), .Y(\u_div/PartRem[53][3] ) );
  CLKINVX1 U244 ( .A(\u_div/PartRem[54][2] ), .Y(\u_div/SumTmp[53][2] ) );
  MXI2X1 U245 ( .A(\u_div/SumTmp[48][2] ), .B(\u_div/PartRem[49][2] ), .S0(
        \u_div/CryTmp[48][6] ), .Y(\u_div/PartRem[48][3] ) );
  CLKINVX1 U246 ( .A(\u_div/PartRem[49][2] ), .Y(\u_div/SumTmp[48][2] ) );
  MXI2X1 U247 ( .A(\u_div/SumTmp[43][2] ), .B(\u_div/PartRem[44][2] ), .S0(
        \u_div/CryTmp[43][6] ), .Y(\u_div/PartRem[43][3] ) );
  CLKINVX1 U248 ( .A(\u_div/PartRem[44][2] ), .Y(\u_div/SumTmp[43][2] ) );
  MXI2X1 U249 ( .A(\u_div/SumTmp[38][2] ), .B(\u_div/PartRem[39][2] ), .S0(
        \u_div/CryTmp[38][6] ), .Y(\u_div/PartRem[38][3] ) );
  CLKINVX1 U250 ( .A(\u_div/PartRem[39][2] ), .Y(\u_div/SumTmp[38][2] ) );
  MXI2X1 U251 ( .A(\u_div/SumTmp[33][2] ), .B(\u_div/PartRem[34][2] ), .S0(
        \u_div/CryTmp[33][6] ), .Y(\u_div/PartRem[33][3] ) );
  CLKINVX1 U252 ( .A(\u_div/PartRem[34][2] ), .Y(\u_div/SumTmp[33][2] ) );
  MXI2X1 U253 ( .A(\u_div/SumTmp[28][2] ), .B(\u_div/PartRem[29][2] ), .S0(
        \u_div/CryTmp[28][6] ), .Y(\u_div/PartRem[28][3] ) );
  CLKINVX1 U254 ( .A(\u_div/PartRem[29][2] ), .Y(\u_div/SumTmp[28][2] ) );
  MXI2X1 U255 ( .A(\u_div/SumTmp[23][2] ), .B(\u_div/PartRem[24][2] ), .S0(
        \u_div/CryTmp[23][6] ), .Y(\u_div/PartRem[23][3] ) );
  CLKINVX1 U256 ( .A(\u_div/PartRem[24][2] ), .Y(\u_div/SumTmp[23][2] ) );
  MXI2X1 U257 ( .A(\u_div/SumTmp[20][2] ), .B(\u_div/PartRem[21][2] ), .S0(
        \u_div/CryTmp[20][6] ), .Y(\u_div/PartRem[20][3] ) );
  CLKINVX1 U258 ( .A(\u_div/PartRem[21][2] ), .Y(\u_div/SumTmp[20][2] ) );
  CLKINVX1 U259 ( .A(\u_div/PartRem[2][2] ), .Y(\u_div/SumTmp[1][2] ) );
  INVX4 U260 ( .A(n2), .Y(n4) );
  INVX4 U261 ( .A(n2), .Y(n5) );
  OR2X2 U262 ( .A(\u_div/PartRem[24][5] ), .B(\u_div/u_add_PartRem_2_23/n2 ), 
        .Y(\u_div/CryTmp[23][6] ) );
  OR2X2 U263 ( .A(\u_div/PartRem[29][5] ), .B(\u_div/u_add_PartRem_2_28/n2 ), 
        .Y(\u_div/CryTmp[28][6] ) );
  OR2X2 U264 ( .A(\u_div/PartRem[34][5] ), .B(\u_div/u_add_PartRem_2_33/n2 ), 
        .Y(\u_div/CryTmp[33][6] ) );
  OR2X2 U265 ( .A(\u_div/PartRem[39][5] ), .B(\u_div/u_add_PartRem_2_38/n2 ), 
        .Y(\u_div/CryTmp[38][6] ) );
  OR2X2 U266 ( .A(\u_div/PartRem[44][5] ), .B(\u_div/u_add_PartRem_2_43/n2 ), 
        .Y(\u_div/CryTmp[43][6] ) );
  OR2X2 U267 ( .A(\u_div/PartRem[49][5] ), .B(\u_div/u_add_PartRem_2_48/n2 ), 
        .Y(\u_div/CryTmp[48][6] ) );
  OR2X2 U268 ( .A(\u_div/PartRem[54][5] ), .B(\u_div/u_add_PartRem_2_53/n2 ), 
        .Y(\u_div/CryTmp[53][6] ) );
  OR2X1 U269 ( .A(\u_div/PartRem[59][5] ), .B(\u_div/u_add_PartRem_2_58/n2 ), 
        .Y(\u_div/CryTmp[58][6] ) );
  XNOR2X1 U270 ( .A(\u_div/PartRem[59][3] ), .B(\u_div/PartRem[59][2] ), .Y(
        \u_div/SumTmp[58][3] ) );
  OR2X1 U271 ( .A(\u_div/PartRem[58][5] ), .B(\u_div/u_add_PartRem_2_57/n2 ), 
        .Y(\u_div/CryTmp[57][6] ) );
  XNOR2X1 U272 ( .A(\u_div/PartRem[58][3] ), .B(\u_div/PartRem[58][2] ), .Y(
        \u_div/SumTmp[57][3] ) );
  OR2X1 U273 ( .A(\u_div/PartRem[57][5] ), .B(\u_div/u_add_PartRem_2_56/n2 ), 
        .Y(\u_div/CryTmp[56][6] ) );
  XNOR2X1 U274 ( .A(\u_div/PartRem[57][3] ), .B(\u_div/PartRem[57][2] ), .Y(
        \u_div/SumTmp[56][3] ) );
  OR2X1 U275 ( .A(\u_div/PartRem[56][5] ), .B(\u_div/u_add_PartRem_2_55/n2 ), 
        .Y(\u_div/CryTmp[55][6] ) );
  XNOR2X1 U276 ( .A(\u_div/PartRem[56][3] ), .B(\u_div/PartRem[56][2] ), .Y(
        \u_div/SumTmp[55][3] ) );
  OR2X1 U277 ( .A(\u_div/PartRem[55][5] ), .B(\u_div/u_add_PartRem_2_54/n2 ), 
        .Y(\u_div/CryTmp[54][6] ) );
  XNOR2X1 U278 ( .A(\u_div/PartRem[55][3] ), .B(\u_div/PartRem[55][2] ), .Y(
        \u_div/SumTmp[54][3] ) );
  XNOR2X1 U279 ( .A(\u_div/PartRem[54][3] ), .B(\u_div/PartRem[54][2] ), .Y(
        \u_div/SumTmp[53][3] ) );
  OR2X1 U280 ( .A(\u_div/PartRem[53][5] ), .B(\u_div/u_add_PartRem_2_52/n2 ), 
        .Y(\u_div/CryTmp[52][6] ) );
  XNOR2X1 U281 ( .A(\u_div/PartRem[53][3] ), .B(\u_div/PartRem[53][2] ), .Y(
        \u_div/SumTmp[52][3] ) );
  XNOR2X1 U282 ( .A(\u_div/PartRem[52][3] ), .B(\u_div/PartRem[52][2] ), .Y(
        \u_div/SumTmp[51][3] ) );
  OR2X1 U283 ( .A(\u_div/PartRem[51][5] ), .B(\u_div/u_add_PartRem_2_50/n2 ), 
        .Y(\u_div/CryTmp[50][6] ) );
  XNOR2X1 U284 ( .A(\u_div/PartRem[51][3] ), .B(\u_div/PartRem[51][2] ), .Y(
        \u_div/SumTmp[50][3] ) );
  OR2X1 U285 ( .A(\u_div/PartRem[51][2] ), .B(\u_div/PartRem[51][3] ), .Y(
        \u_div/u_add_PartRem_2_50/n3 ) );
  OR2X1 U286 ( .A(\u_div/PartRem[50][5] ), .B(\u_div/u_add_PartRem_2_49/n2 ), 
        .Y(\u_div/CryTmp[49][6] ) );
  XNOR2X1 U287 ( .A(\u_div/PartRem[50][3] ), .B(\u_div/PartRem[50][2] ), .Y(
        \u_div/SumTmp[49][3] ) );
  XNOR2X1 U288 ( .A(\u_div/PartRem[49][3] ), .B(\u_div/PartRem[49][2] ), .Y(
        \u_div/SumTmp[48][3] ) );
  OR2X1 U289 ( .A(\u_div/PartRem[48][5] ), .B(\u_div/u_add_PartRem_2_47/n2 ), 
        .Y(\u_div/CryTmp[47][6] ) );
  XNOR2X1 U290 ( .A(\u_div/PartRem[48][3] ), .B(\u_div/PartRem[48][2] ), .Y(
        \u_div/SumTmp[47][3] ) );
  XNOR2X1 U291 ( .A(\u_div/PartRem[47][3] ), .B(\u_div/PartRem[47][2] ), .Y(
        \u_div/SumTmp[46][3] ) );
  OR2X1 U292 ( .A(\u_div/PartRem[46][5] ), .B(\u_div/u_add_PartRem_2_45/n2 ), 
        .Y(\u_div/CryTmp[45][6] ) );
  XNOR2X1 U293 ( .A(\u_div/PartRem[46][3] ), .B(\u_div/PartRem[46][2] ), .Y(
        \u_div/SumTmp[45][3] ) );
  OR2X1 U294 ( .A(\u_div/PartRem[46][2] ), .B(\u_div/PartRem[46][3] ), .Y(
        \u_div/u_add_PartRem_2_45/n3 ) );
  OR2X1 U295 ( .A(\u_div/PartRem[45][5] ), .B(\u_div/u_add_PartRem_2_44/n2 ), 
        .Y(\u_div/CryTmp[44][6] ) );
  XNOR2X1 U296 ( .A(\u_div/PartRem[45][3] ), .B(\u_div/PartRem[45][2] ), .Y(
        \u_div/SumTmp[44][3] ) );
  XNOR2X1 U297 ( .A(\u_div/PartRem[44][3] ), .B(\u_div/PartRem[44][2] ), .Y(
        \u_div/SumTmp[43][3] ) );
  OR2X1 U298 ( .A(\u_div/PartRem[43][5] ), .B(\u_div/u_add_PartRem_2_42/n2 ), 
        .Y(\u_div/CryTmp[42][6] ) );
  XNOR2X1 U299 ( .A(\u_div/PartRem[43][3] ), .B(\u_div/PartRem[43][2] ), .Y(
        \u_div/SumTmp[42][3] ) );
  OR2X1 U300 ( .A(\u_div/PartRem[42][5] ), .B(\u_div/u_add_PartRem_2_41/n2 ), 
        .Y(\u_div/CryTmp[41][6] ) );
  XNOR2X1 U301 ( .A(\u_div/PartRem[42][3] ), .B(\u_div/PartRem[42][2] ), .Y(
        \u_div/SumTmp[41][3] ) );
  OR2X1 U302 ( .A(\u_div/PartRem[41][5] ), .B(\u_div/u_add_PartRem_2_40/n2 ), 
        .Y(\u_div/CryTmp[40][6] ) );
  XNOR2X1 U303 ( .A(\u_div/PartRem[41][3] ), .B(\u_div/PartRem[41][2] ), .Y(
        \u_div/SumTmp[40][3] ) );
  OR2X1 U304 ( .A(\u_div/PartRem[41][2] ), .B(\u_div/PartRem[41][3] ), .Y(
        \u_div/u_add_PartRem_2_40/n3 ) );
  OR2X1 U305 ( .A(\u_div/PartRem[40][5] ), .B(\u_div/u_add_PartRem_2_39/n2 ), 
        .Y(\u_div/CryTmp[39][6] ) );
  XNOR2X1 U306 ( .A(\u_div/PartRem[40][3] ), .B(\u_div/PartRem[40][2] ), .Y(
        \u_div/SumTmp[39][3] ) );
  XNOR2X1 U307 ( .A(\u_div/PartRem[39][3] ), .B(\u_div/PartRem[39][2] ), .Y(
        \u_div/SumTmp[38][3] ) );
  OR2X1 U308 ( .A(\u_div/PartRem[38][5] ), .B(\u_div/u_add_PartRem_2_37/n2 ), 
        .Y(\u_div/CryTmp[37][6] ) );
  XNOR2X1 U309 ( .A(\u_div/PartRem[38][3] ), .B(\u_div/PartRem[38][2] ), .Y(
        \u_div/SumTmp[37][3] ) );
  XNOR2X1 U310 ( .A(\u_div/PartRem[37][3] ), .B(\u_div/PartRem[37][2] ), .Y(
        \u_div/SumTmp[36][3] ) );
  OR2X1 U311 ( .A(\u_div/PartRem[36][5] ), .B(\u_div/u_add_PartRem_2_35/n2 ), 
        .Y(\u_div/CryTmp[35][6] ) );
  XNOR2X1 U312 ( .A(\u_div/PartRem[36][3] ), .B(\u_div/PartRem[36][2] ), .Y(
        \u_div/SumTmp[35][3] ) );
  OR2X1 U313 ( .A(\u_div/PartRem[36][2] ), .B(\u_div/PartRem[36][3] ), .Y(
        \u_div/u_add_PartRem_2_35/n3 ) );
  OR2X1 U314 ( .A(\u_div/PartRem[35][5] ), .B(\u_div/u_add_PartRem_2_34/n2 ), 
        .Y(\u_div/CryTmp[34][6] ) );
  XNOR2X1 U315 ( .A(\u_div/PartRem[35][3] ), .B(\u_div/PartRem[35][2] ), .Y(
        \u_div/SumTmp[34][3] ) );
  XNOR2X1 U316 ( .A(\u_div/PartRem[34][3] ), .B(\u_div/PartRem[34][2] ), .Y(
        \u_div/SumTmp[33][3] ) );
  OR2X1 U317 ( .A(\u_div/PartRem[33][5] ), .B(\u_div/u_add_PartRem_2_32/n2 ), 
        .Y(\u_div/CryTmp[32][6] ) );
  XNOR2X1 U318 ( .A(\u_div/PartRem[33][3] ), .B(\u_div/PartRem[33][2] ), .Y(
        \u_div/SumTmp[32][3] ) );
  OR2X1 U319 ( .A(\u_div/PartRem[32][5] ), .B(\u_div/u_add_PartRem_2_31/n2 ), 
        .Y(\u_div/CryTmp[31][6] ) );
  XNOR2X1 U320 ( .A(\u_div/PartRem[32][3] ), .B(\u_div/PartRem[32][2] ), .Y(
        \u_div/SumTmp[31][3] ) );
  OR2X1 U321 ( .A(\u_div/PartRem[31][5] ), .B(\u_div/u_add_PartRem_2_30/n2 ), 
        .Y(\u_div/CryTmp[30][6] ) );
  XNOR2X1 U322 ( .A(\u_div/PartRem[31][3] ), .B(\u_div/PartRem[31][2] ), .Y(
        \u_div/SumTmp[30][3] ) );
  OR2X1 U323 ( .A(\u_div/PartRem[31][2] ), .B(\u_div/PartRem[31][3] ), .Y(
        \u_div/u_add_PartRem_2_30/n3 ) );
  OR2X1 U324 ( .A(\u_div/PartRem[30][5] ), .B(\u_div/u_add_PartRem_2_29/n2 ), 
        .Y(\u_div/CryTmp[29][6] ) );
  XNOR2X1 U325 ( .A(\u_div/PartRem[30][3] ), .B(\u_div/PartRem[30][2] ), .Y(
        \u_div/SumTmp[29][3] ) );
  XNOR2X1 U326 ( .A(\u_div/PartRem[29][3] ), .B(\u_div/PartRem[29][2] ), .Y(
        \u_div/SumTmp[28][3] ) );
  OR2X1 U327 ( .A(\u_div/PartRem[28][5] ), .B(\u_div/u_add_PartRem_2_27/n2 ), 
        .Y(\u_div/CryTmp[27][6] ) );
  XNOR2X1 U328 ( .A(\u_div/PartRem[28][3] ), .B(\u_div/PartRem[28][2] ), .Y(
        \u_div/SumTmp[27][3] ) );
  XNOR2X1 U329 ( .A(\u_div/PartRem[27][3] ), .B(\u_div/PartRem[27][2] ), .Y(
        \u_div/SumTmp[26][3] ) );
  OR2X1 U330 ( .A(\u_div/PartRem[26][5] ), .B(\u_div/u_add_PartRem_2_25/n2 ), 
        .Y(\u_div/CryTmp[25][6] ) );
  XNOR2X1 U331 ( .A(\u_div/PartRem[26][3] ), .B(\u_div/PartRem[26][2] ), .Y(
        \u_div/SumTmp[25][3] ) );
  OR2X1 U332 ( .A(\u_div/PartRem[26][2] ), .B(\u_div/PartRem[26][3] ), .Y(
        \u_div/u_add_PartRem_2_25/n3 ) );
  OR2X1 U333 ( .A(\u_div/PartRem[25][5] ), .B(\u_div/u_add_PartRem_2_24/n2 ), 
        .Y(\u_div/CryTmp[24][6] ) );
  XNOR2X1 U334 ( .A(\u_div/PartRem[25][3] ), .B(\u_div/PartRem[25][2] ), .Y(
        \u_div/SumTmp[24][3] ) );
  XNOR2X1 U335 ( .A(\u_div/PartRem[24][3] ), .B(\u_div/PartRem[24][2] ), .Y(
        \u_div/SumTmp[23][3] ) );
  OR2X1 U336 ( .A(\u_div/PartRem[23][5] ), .B(\u_div/u_add_PartRem_2_22/n2 ), 
        .Y(\u_div/CryTmp[22][6] ) );
  XNOR2X1 U337 ( .A(\u_div/PartRem[23][3] ), .B(\u_div/PartRem[23][2] ), .Y(
        \u_div/SumTmp[22][3] ) );
  OR2X1 U338 ( .A(\u_div/PartRem[22][5] ), .B(\u_div/u_add_PartRem_2_21/n2 ), 
        .Y(\u_div/CryTmp[21][6] ) );
  XNOR2X1 U339 ( .A(\u_div/PartRem[22][3] ), .B(\u_div/PartRem[22][2] ), .Y(
        \u_div/SumTmp[21][3] ) );
  XNOR2X1 U340 ( .A(\u_div/PartRem[21][3] ), .B(\u_div/PartRem[21][2] ), .Y(
        \u_div/SumTmp[20][3] ) );
  OR2X1 U341 ( .A(\u_div/PartRem[20][5] ), .B(\u_div/u_add_PartRem_2_19/n2 ), 
        .Y(\u_div/CryTmp[19][6] ) );
  XNOR2X1 U342 ( .A(\u_div/PartRem[20][3] ), .B(\u_div/PartRem[20][2] ), .Y(
        \u_div/SumTmp[19][3] ) );
  XNOR2X1 U343 ( .A(\u_div/PartRem[19][3] ), .B(\u_div/PartRem[19][2] ), .Y(
        \u_div/SumTmp[18][3] ) );
  OR2X1 U344 ( .A(\u_div/PartRem[18][5] ), .B(\u_div/u_add_PartRem_2_17/n2 ), 
        .Y(\u_div/CryTmp[17][6] ) );
  XNOR2X1 U345 ( .A(\u_div/PartRem[18][3] ), .B(\u_div/PartRem[18][2] ), .Y(
        \u_div/SumTmp[17][3] ) );
  OR2X1 U346 ( .A(\u_div/PartRem[17][5] ), .B(\u_div/u_add_PartRem_2_16/n2 ), 
        .Y(\u_div/CryTmp[16][6] ) );
  XNOR2X1 U347 ( .A(\u_div/PartRem[17][3] ), .B(\u_div/PartRem[17][2] ), .Y(
        \u_div/SumTmp[16][3] ) );
  OR2X1 U348 ( .A(\u_div/PartRem[16][5] ), .B(\u_div/u_add_PartRem_2_15/n2 ), 
        .Y(\u_div/CryTmp[15][6] ) );
  XNOR2X1 U349 ( .A(\u_div/PartRem[16][3] ), .B(\u_div/PartRem[16][2] ), .Y(
        \u_div/SumTmp[15][3] ) );
  OR2X1 U350 ( .A(\u_div/PartRem[15][5] ), .B(\u_div/u_add_PartRem_2_14/n2 ), 
        .Y(\u_div/CryTmp[14][6] ) );
  XNOR2X1 U351 ( .A(\u_div/PartRem[15][3] ), .B(\u_div/PartRem[15][2] ), .Y(
        \u_div/SumTmp[14][3] ) );
  XNOR2X1 U352 ( .A(\u_div/PartRem[14][3] ), .B(\u_div/PartRem[14][2] ), .Y(
        \u_div/SumTmp[13][3] ) );
  OR2X1 U353 ( .A(\u_div/PartRem[13][5] ), .B(\u_div/u_add_PartRem_2_12/n2 ), 
        .Y(\u_div/CryTmp[12][6] ) );
  XNOR2X1 U354 ( .A(\u_div/PartRem[13][3] ), .B(\u_div/PartRem[13][2] ), .Y(
        \u_div/SumTmp[12][3] ) );
  OR2X1 U355 ( .A(\u_div/PartRem[12][5] ), .B(\u_div/u_add_PartRem_2_11/n2 ), 
        .Y(\u_div/CryTmp[11][6] ) );
  XNOR2X1 U356 ( .A(\u_div/PartRem[12][3] ), .B(\u_div/PartRem[12][2] ), .Y(
        \u_div/SumTmp[11][3] ) );
  OR2X1 U357 ( .A(\u_div/PartRem[11][5] ), .B(\u_div/u_add_PartRem_2_10/n2 ), 
        .Y(\u_div/CryTmp[10][6] ) );
  XNOR2X1 U358 ( .A(\u_div/PartRem[11][3] ), .B(\u_div/PartRem[11][2] ), .Y(
        \u_div/SumTmp[10][3] ) );
  OR2X1 U359 ( .A(\u_div/PartRem[10][5] ), .B(\u_div/u_add_PartRem_2_9/n2 ), 
        .Y(\u_div/CryTmp[9][6] ) );
  XNOR2X1 U360 ( .A(\u_div/PartRem[10][3] ), .B(\u_div/PartRem[10][2] ), .Y(
        \u_div/SumTmp[9][3] ) );
  XNOR2X1 U361 ( .A(\u_div/PartRem[9][3] ), .B(\u_div/PartRem[9][2] ), .Y(
        \u_div/SumTmp[8][3] ) );
  XNOR2X1 U362 ( .A(\u_div/PartRem[8][3] ), .B(\u_div/PartRem[8][2] ), .Y(
        \u_div/SumTmp[7][3] ) );
  OR2X1 U363 ( .A(\u_div/PartRem[7][5] ), .B(\u_div/u_add_PartRem_2_6/n2 ), 
        .Y(\u_div/CryTmp[6][6] ) );
  XNOR2X1 U364 ( .A(\u_div/PartRem[7][3] ), .B(\u_div/PartRem[7][2] ), .Y(
        \u_div/SumTmp[6][3] ) );
  OR2X1 U365 ( .A(\u_div/PartRem[6][5] ), .B(\u_div/u_add_PartRem_2_5/n2 ), 
        .Y(\u_div/CryTmp[5][6] ) );
  XNOR2X1 U366 ( .A(\u_div/PartRem[6][3] ), .B(\u_div/PartRem[6][2] ), .Y(
        \u_div/SumTmp[5][3] ) );
  XNOR2X1 U367 ( .A(\u_div/PartRem[5][3] ), .B(\u_div/PartRem[5][2] ), .Y(
        \u_div/SumTmp[4][3] ) );
  OR2X1 U368 ( .A(\u_div/PartRem[4][5] ), .B(\u_div/u_add_PartRem_2_3/n2 ), 
        .Y(\u_div/CryTmp[3][6] ) );
  XNOR2X1 U369 ( .A(\u_div/PartRem[4][3] ), .B(\u_div/PartRem[4][2] ), .Y(
        \u_div/SumTmp[3][3] ) );
  OR2X1 U370 ( .A(\u_div/PartRem[4][2] ), .B(\u_div/PartRem[4][3] ), .Y(
        \u_div/u_add_PartRem_2_3/n3 ) );
  XNOR2X1 U371 ( .A(\u_div/PartRem[3][3] ), .B(\u_div/PartRem[3][2] ), .Y(
        \u_div/SumTmp[2][3] ) );
  XNOR2X1 U372 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/PartRem[2][2] ), .Y(
        \u_div/SumTmp[1][3] ) );
  XNOR2X1 U373 ( .A(\u_div/PartRem[63][0] ), .B(\u_div/PartRem[62][0] ), .Y(
        \u_div/SumTmp[59][3] ) );
  XOR2X1 U374 ( .A(\u_div/CryTmp[9][6] ), .B(n3), .Y(\u_div/QInv[9] ) );
  XOR2X1 U375 ( .A(\u_div/CryTmp[7][6] ), .B(n4), .Y(\u_div/QInv[7] ) );
  XOR2X1 U376 ( .A(\u_div/CryTmp[59][6] ), .B(n3), .Y(\u_div/QInv[59] ) );
  XOR2X1 U377 ( .A(\u_div/CryTmp[58][6] ), .B(n5), .Y(\u_div/QInv[58] ) );
  XOR2X1 U378 ( .A(\u_div/CryTmp[57][6] ), .B(n4), .Y(\u_div/QInv[57] ) );
  XOR2X1 U379 ( .A(\u_div/CryTmp[56][6] ), .B(n3), .Y(\u_div/QInv[56] ) );
  XOR2X1 U380 ( .A(\u_div/CryTmp[54][6] ), .B(n4), .Y(\u_div/QInv[54] ) );
  XOR2X1 U381 ( .A(\u_div/CryTmp[53][6] ), .B(n3), .Y(\u_div/QInv[53] ) );
  XOR2X1 U382 ( .A(\u_div/CryTmp[52][6] ), .B(n5), .Y(\u_div/QInv[52] ) );
  XOR2X1 U383 ( .A(\u_div/CryTmp[49][6] ), .B(n4), .Y(\u_div/QInv[49] ) );
  XOR2X1 U384 ( .A(\u_div/CryTmp[48][6] ), .B(n3), .Y(\u_div/QInv[48] ) );
  XOR2X1 U385 ( .A(\u_div/CryTmp[47][6] ), .B(n5), .Y(\u_div/QInv[47] ) );
  XOR2X1 U386 ( .A(\u_div/CryTmp[46][6] ), .B(n4), .Y(\u_div/QInv[46] ) );
  XOR2X1 U387 ( .A(\u_div/CryTmp[45][6] ), .B(n3), .Y(\u_div/QInv[45] ) );
  XOR2X1 U388 ( .A(\u_div/CryTmp[39][6] ), .B(n5), .Y(\u_div/QInv[39] ) );
  XOR2X1 U389 ( .A(\u_div/CryTmp[38][6] ), .B(n4), .Y(\u_div/QInv[38] ) );
  XOR2X1 U390 ( .A(\u_div/CryTmp[37][6] ), .B(n3), .Y(\u_div/QInv[37] ) );
  XOR2X1 U391 ( .A(\u_div/CryTmp[36][6] ), .B(n5), .Y(\u_div/QInv[36] ) );
  XOR2X1 U392 ( .A(\u_div/CryTmp[35][6] ), .B(n4), .Y(\u_div/QInv[35] ) );
  XOR2X1 U393 ( .A(\u_div/CryTmp[34][6] ), .B(n5), .Y(\u_div/QInv[34] ) );
  XOR2X1 U394 ( .A(\u_div/CryTmp[33][6] ), .B(n4), .Y(\u_div/QInv[33] ) );
  XOR2X1 U395 ( .A(\u_div/CryTmp[32][6] ), .B(n3), .Y(\u_div/QInv[32] ) );
  XOR2X1 U396 ( .A(\u_div/CryTmp[29][6] ), .B(n5), .Y(\u_div/QInv[29] ) );
  XOR2X1 U397 ( .A(\u_div/CryTmp[28][6] ), .B(n4), .Y(\u_div/QInv[28] ) );
  XOR2X1 U398 ( .A(\u_div/CryTmp[27][6] ), .B(n3), .Y(\u_div/QInv[27] ) );
  XOR2X1 U399 ( .A(\u_div/CryTmp[26][6] ), .B(n5), .Y(\u_div/QInv[26] ) );
  XOR2X1 U400 ( .A(\u_div/CryTmp[25][6] ), .B(n4), .Y(\u_div/QInv[25] ) );
  XOR2X1 U401 ( .A(\u_div/CryTmp[24][6] ), .B(n3), .Y(\u_div/QInv[24] ) );
  XOR2X1 U402 ( .A(\u_div/CryTmp[23][6] ), .B(n5), .Y(\u_div/QInv[23] ) );
  XOR2X1 U403 ( .A(\u_div/CryTmp[22][6] ), .B(n4), .Y(\u_div/QInv[22] ) );
  XOR2X1 U404 ( .A(\u_div/CryTmp[1][6] ), .B(n4), .Y(\u_div/QInv[1] ) );
  XOR2X1 U405 ( .A(\u_div/CryTmp[19][6] ), .B(n3), .Y(\u_div/QInv[19] ) );
  XOR2X1 U406 ( .A(\u_div/CryTmp[18][6] ), .B(n5), .Y(\u_div/QInv[18] ) );
  XOR2X1 U407 ( .A(\u_div/CryTmp[17][6] ), .B(n4), .Y(\u_div/QInv[17] ) );
  XOR2X1 U408 ( .A(\u_div/CryTmp[15][6] ), .B(n4), .Y(\u_div/QInv[15] ) );
  XOR2X1 U409 ( .A(\u_div/CryTmp[14][6] ), .B(n5), .Y(\u_div/QInv[14] ) );
endmodule


module GSIM_DW01_inc_6 ( A, SUM );
  input [63:0] A;
  output [63:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;

  NOR3BX1 U2 ( .AN(A[15]), .B(n12), .C(n72), .Y(n70) );
  NOR3BX1 U3 ( .AN(A[19]), .B(n11), .C(n68), .Y(n66) );
  NOR3BX1 U4 ( .AN(A[23]), .B(n10), .C(n64), .Y(n62) );
  NOR3BX1 U5 ( .AN(A[11]), .B(n13), .C(n76), .Y(n74) );
  NOR3BX1 U6 ( .AN(A[7]), .B(n14), .C(n19), .Y(n17) );
  NOR3BX1 U7 ( .AN(A[27]), .B(n9), .C(n60), .Y(n58) );
  NOR3BX1 U8 ( .AN(A[31]), .B(n8), .C(n56), .Y(n54) );
  NOR3BX1 U9 ( .AN(A[35]), .B(n7), .C(n52), .Y(n50) );
  NOR3BX1 U10 ( .AN(A[39]), .B(n6), .C(n46), .Y(n44) );
  NOR3BX1 U11 ( .AN(A[43]), .B(n5), .C(n42), .Y(n40) );
  NOR3BX1 U12 ( .AN(A[47]), .B(n4), .C(n38), .Y(n36) );
  NOR3BX1 U13 ( .AN(A[51]), .B(n3), .C(n34), .Y(n32) );
  NOR3BX1 U14 ( .AN(A[55]), .B(n2), .C(n30), .Y(n28) );
  NOR3BX1 U15 ( .AN(A[59]), .B(n1), .C(n24), .Y(n22) );
  NAND2XL U16 ( .A(A[60]), .B(n22), .Y(n23) );
  NAND3X1 U17 ( .A(A[4]), .B(n26), .C(A[5]), .Y(n19) );
  NOR3BX1 U18 ( .AN(A[3]), .B(n15), .C(n48), .Y(n26) );
  NOR2XL U19 ( .A(n24), .B(n1), .Y(n27) );
  NAND2XL U20 ( .A(A[56]), .B(n28), .Y(n29) );
  NOR2XL U21 ( .A(n30), .B(n2), .Y(n31) );
  NAND2XL U22 ( .A(A[52]), .B(n32), .Y(n33) );
  NOR2XL U23 ( .A(n34), .B(n3), .Y(n35) );
  NAND2XL U24 ( .A(A[48]), .B(n36), .Y(n37) );
  NOR2XL U25 ( .A(n38), .B(n4), .Y(n39) );
  NAND2XL U26 ( .A(A[44]), .B(n40), .Y(n41) );
  NOR2XL U27 ( .A(n42), .B(n5), .Y(n43) );
  NAND2XL U28 ( .A(A[40]), .B(n44), .Y(n45) );
  NOR2XL U29 ( .A(n46), .B(n6), .Y(n49) );
  NAND2XL U30 ( .A(A[36]), .B(n50), .Y(n51) );
  NOR2XL U31 ( .A(n52), .B(n7), .Y(n53) );
  NAND2XL U32 ( .A(A[32]), .B(n54), .Y(n55) );
  NOR2XL U33 ( .A(n56), .B(n8), .Y(n57) );
  NAND2XL U34 ( .A(A[28]), .B(n58), .Y(n59) );
  NOR2XL U35 ( .A(n60), .B(n9), .Y(n61) );
  NAND2XL U36 ( .A(A[24]), .B(n62), .Y(n63) );
  NOR2XL U37 ( .A(n64), .B(n10), .Y(n65) );
  NAND2XL U38 ( .A(A[20]), .B(n66), .Y(n67) );
  NOR2XL U39 ( .A(n68), .B(n11), .Y(n69) );
  NAND2XL U40 ( .A(A[16]), .B(n70), .Y(n71) );
  NOR2XL U41 ( .A(n72), .B(n12), .Y(n73) );
  NAND2XL U42 ( .A(A[12]), .B(n74), .Y(n75) );
  NOR2XL U43 ( .A(n76), .B(n13), .Y(n77) );
  NAND2XL U44 ( .A(A[8]), .B(n17), .Y(n16) );
  NOR2XL U45 ( .A(n19), .B(n14), .Y(n18) );
  NAND2XL U46 ( .A(A[4]), .B(n26), .Y(n25) );
  XOR2XL U47 ( .A(A[60]), .B(n22), .Y(SUM[60]) );
  XNOR2XL U48 ( .A(A[61]), .B(n23), .Y(SUM[61]) );
  XNOR2XL U49 ( .A(A[62]), .B(n21), .Y(SUM[62]) );
  NOR2XL U50 ( .A(n48), .B(n15), .Y(n47) );
  CLKINVX1 U51 ( .A(A[58]), .Y(n1) );
  CLKINVX1 U52 ( .A(A[42]), .Y(n5) );
  CLKINVX1 U53 ( .A(A[46]), .Y(n4) );
  CLKINVX1 U54 ( .A(A[54]), .Y(n2) );
  CLKINVX1 U55 ( .A(A[38]), .Y(n6) );
  CLKINVX1 U56 ( .A(A[34]), .Y(n7) );
  CLKINVX1 U57 ( .A(A[30]), .Y(n8) );
  CLKINVX1 U58 ( .A(A[26]), .Y(n9) );
  CLKINVX1 U59 ( .A(A[22]), .Y(n10) );
  CLKINVX1 U60 ( .A(A[18]), .Y(n11) );
  CLKINVX1 U61 ( .A(A[14]), .Y(n12) );
  CLKINVX1 U62 ( .A(A[2]), .Y(n15) );
  CLKINVX1 U63 ( .A(A[50]), .Y(n3) );
  CLKINVX1 U64 ( .A(A[10]), .Y(n13) );
  CLKINVX1 U65 ( .A(A[6]), .Y(n14) );
  XNOR2X1 U66 ( .A(A[9]), .B(n16), .Y(SUM[9]) );
  XOR2X1 U67 ( .A(A[8]), .B(n17), .Y(SUM[8]) );
  XOR2X1 U68 ( .A(A[7]), .B(n18), .Y(SUM[7]) );
  XOR2X1 U69 ( .A(n14), .B(n19), .Y(SUM[6]) );
  XOR2X1 U70 ( .A(A[63]), .B(n20), .Y(SUM[63]) );
  NOR2BX1 U71 ( .AN(A[62]), .B(n21), .Y(n20) );
  NAND3X1 U72 ( .A(A[60]), .B(n22), .C(A[61]), .Y(n21) );
  XNOR2X1 U73 ( .A(A[5]), .B(n25), .Y(SUM[5]) );
  XOR2X1 U74 ( .A(A[59]), .B(n27), .Y(SUM[59]) );
  XOR2X1 U75 ( .A(n1), .B(n24), .Y(SUM[58]) );
  NAND3X1 U76 ( .A(A[56]), .B(n28), .C(A[57]), .Y(n24) );
  XNOR2X1 U77 ( .A(A[57]), .B(n29), .Y(SUM[57]) );
  XOR2X1 U78 ( .A(A[56]), .B(n28), .Y(SUM[56]) );
  XOR2X1 U79 ( .A(A[55]), .B(n31), .Y(SUM[55]) );
  XOR2X1 U80 ( .A(n2), .B(n30), .Y(SUM[54]) );
  NAND3X1 U81 ( .A(A[52]), .B(n32), .C(A[53]), .Y(n30) );
  XNOR2X1 U82 ( .A(A[53]), .B(n33), .Y(SUM[53]) );
  XOR2X1 U83 ( .A(A[52]), .B(n32), .Y(SUM[52]) );
  XOR2X1 U84 ( .A(A[51]), .B(n35), .Y(SUM[51]) );
  XOR2X1 U85 ( .A(n3), .B(n34), .Y(SUM[50]) );
  NAND3X1 U86 ( .A(A[48]), .B(n36), .C(A[49]), .Y(n34) );
  XOR2X1 U87 ( .A(A[4]), .B(n26), .Y(SUM[4]) );
  XNOR2X1 U88 ( .A(A[49]), .B(n37), .Y(SUM[49]) );
  XOR2X1 U89 ( .A(A[48]), .B(n36), .Y(SUM[48]) );
  XOR2X1 U90 ( .A(A[47]), .B(n39), .Y(SUM[47]) );
  XOR2X1 U91 ( .A(n4), .B(n38), .Y(SUM[46]) );
  NAND3X1 U92 ( .A(A[44]), .B(n40), .C(A[45]), .Y(n38) );
  XNOR2X1 U93 ( .A(A[45]), .B(n41), .Y(SUM[45]) );
  XOR2X1 U94 ( .A(A[44]), .B(n40), .Y(SUM[44]) );
  XOR2X1 U95 ( .A(A[43]), .B(n43), .Y(SUM[43]) );
  XOR2X1 U96 ( .A(n5), .B(n42), .Y(SUM[42]) );
  NAND3X1 U97 ( .A(A[40]), .B(n44), .C(A[41]), .Y(n42) );
  XNOR2X1 U98 ( .A(A[41]), .B(n45), .Y(SUM[41]) );
  XOR2X1 U99 ( .A(A[40]), .B(n44), .Y(SUM[40]) );
  XOR2X1 U100 ( .A(A[3]), .B(n47), .Y(SUM[3]) );
  XOR2X1 U101 ( .A(A[39]), .B(n49), .Y(SUM[39]) );
  XOR2X1 U102 ( .A(n6), .B(n46), .Y(SUM[38]) );
  NAND3X1 U103 ( .A(A[36]), .B(n50), .C(A[37]), .Y(n46) );
  XNOR2X1 U104 ( .A(A[37]), .B(n51), .Y(SUM[37]) );
  XOR2X1 U105 ( .A(A[36]), .B(n50), .Y(SUM[36]) );
  XOR2X1 U106 ( .A(A[35]), .B(n53), .Y(SUM[35]) );
  XOR2X1 U107 ( .A(n7), .B(n52), .Y(SUM[34]) );
  NAND3X1 U108 ( .A(A[32]), .B(n54), .C(A[33]), .Y(n52) );
  XNOR2X1 U109 ( .A(A[33]), .B(n55), .Y(SUM[33]) );
  XOR2X1 U110 ( .A(A[32]), .B(n54), .Y(SUM[32]) );
  XOR2X1 U111 ( .A(A[31]), .B(n57), .Y(SUM[31]) );
  XOR2X1 U112 ( .A(n8), .B(n56), .Y(SUM[30]) );
  NAND3X1 U113 ( .A(A[28]), .B(n58), .C(A[29]), .Y(n56) );
  XOR2X1 U114 ( .A(n15), .B(n48), .Y(SUM[2]) );
  XNOR2X1 U115 ( .A(A[29]), .B(n59), .Y(SUM[29]) );
  XOR2X1 U116 ( .A(A[28]), .B(n58), .Y(SUM[28]) );
  XOR2X1 U117 ( .A(A[27]), .B(n61), .Y(SUM[27]) );
  XOR2X1 U118 ( .A(n9), .B(n60), .Y(SUM[26]) );
  NAND3X1 U119 ( .A(A[24]), .B(n62), .C(A[25]), .Y(n60) );
  XNOR2X1 U120 ( .A(A[25]), .B(n63), .Y(SUM[25]) );
  XOR2X1 U121 ( .A(A[24]), .B(n62), .Y(SUM[24]) );
  XOR2X1 U122 ( .A(A[23]), .B(n65), .Y(SUM[23]) );
  XOR2X1 U123 ( .A(n10), .B(n64), .Y(SUM[22]) );
  NAND3X1 U124 ( .A(A[20]), .B(n66), .C(A[21]), .Y(n64) );
  XNOR2X1 U125 ( .A(A[21]), .B(n67), .Y(SUM[21]) );
  XOR2X1 U126 ( .A(A[20]), .B(n66), .Y(SUM[20]) );
  XOR2X1 U127 ( .A(A[19]), .B(n69), .Y(SUM[19]) );
  XOR2X1 U128 ( .A(n11), .B(n68), .Y(SUM[18]) );
  NAND3X1 U129 ( .A(A[16]), .B(n70), .C(A[17]), .Y(n68) );
  XNOR2X1 U130 ( .A(A[17]), .B(n71), .Y(SUM[17]) );
  XOR2X1 U131 ( .A(A[16]), .B(n70), .Y(SUM[16]) );
  XOR2X1 U132 ( .A(A[15]), .B(n73), .Y(SUM[15]) );
  XOR2X1 U133 ( .A(n12), .B(n72), .Y(SUM[14]) );
  NAND3X1 U134 ( .A(A[12]), .B(n74), .C(A[13]), .Y(n72) );
  XNOR2X1 U135 ( .A(A[13]), .B(n75), .Y(SUM[13]) );
  XOR2X1 U136 ( .A(A[12]), .B(n74), .Y(SUM[12]) );
  XOR2X1 U137 ( .A(A[11]), .B(n77), .Y(SUM[11]) );
  XOR2X1 U138 ( .A(n13), .B(n76), .Y(SUM[10]) );
  NAND3X1 U139 ( .A(A[8]), .B(n17), .C(A[9]), .Y(n76) );
  NAND2X1 U140 ( .A(A[1]), .B(A[0]), .Y(n48) );
endmodule


module GSIM_DW01_absval_4 ( A, ABSVAL );
  input [63:0] A;
  output [63:0] ABSVAL;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68;
  wire   [63:0] AMUX1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  GSIM_DW01_inc_6 NEG ( .A({n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
        n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
        n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
        n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
        n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68}), .SUM({
        AMUX1[63:2], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1}) );
  CLKINVX1 U1 ( .A(A[61]), .Y(n7) );
  CLKMX2X2 U2 ( .A(A[61]), .B(AMUX1[61]), .S0(n4), .Y(ABSVAL[61]) );
  INVX3 U3 ( .A(n5), .Y(n4) );
  INVX3 U4 ( .A(n5), .Y(n3) );
  INVX3 U5 ( .A(n5), .Y(n2) );
  INVX3 U6 ( .A(n5), .Y(n1) );
  CLKINVX1 U7 ( .A(A[63]), .Y(n5) );
  CLKINVX1 U8 ( .A(A[58]), .Y(n10) );
  CLKINVX1 U9 ( .A(A[42]), .Y(n26) );
  CLKINVX1 U10 ( .A(A[45]), .Y(n23) );
  CLKINVX1 U11 ( .A(A[62]), .Y(n6) );
  CLKINVX1 U12 ( .A(A[59]), .Y(n9) );
  CLKINVX1 U13 ( .A(A[55]), .Y(n13) );
  CLKINVX1 U14 ( .A(A[51]), .Y(n17) );
  CLKINVX1 U15 ( .A(A[47]), .Y(n21) );
  CLKINVX1 U16 ( .A(A[43]), .Y(n25) );
  CLKINVX1 U17 ( .A(A[39]), .Y(n29) );
  CLKINVX1 U18 ( .A(A[35]), .Y(n33) );
  CLKINVX1 U19 ( .A(A[31]), .Y(n37) );
  CLKINVX1 U20 ( .A(A[27]), .Y(n41) );
  CLKINVX1 U21 ( .A(A[46]), .Y(n22) );
  CLKINVX1 U22 ( .A(A[60]), .Y(n8) );
  CLKINVX1 U23 ( .A(A[56]), .Y(n12) );
  CLKINVX1 U24 ( .A(A[52]), .Y(n16) );
  CLKINVX1 U25 ( .A(A[48]), .Y(n20) );
  CLKINVX1 U26 ( .A(A[44]), .Y(n24) );
  CLKINVX1 U27 ( .A(A[40]), .Y(n28) );
  CLKINVX1 U28 ( .A(A[36]), .Y(n32) );
  CLKINVX1 U29 ( .A(A[32]), .Y(n36) );
  CLKINVX1 U30 ( .A(A[28]), .Y(n40) );
  CLKINVX1 U31 ( .A(A[54]), .Y(n14) );
  CLKINVX1 U32 ( .A(A[38]), .Y(n30) );
  CLKINVX1 U33 ( .A(A[34]), .Y(n34) );
  CLKINVX1 U34 ( .A(A[30]), .Y(n38) );
  CLKINVX1 U35 ( .A(A[26]), .Y(n42) );
  CLKINVX1 U36 ( .A(A[22]), .Y(n46) );
  CLKINVX1 U37 ( .A(A[18]), .Y(n50) );
  CLKINVX1 U38 ( .A(A[14]), .Y(n54) );
  CLKINVX1 U39 ( .A(A[2]), .Y(n66) );
  CLKINVX1 U40 ( .A(A[57]), .Y(n11) );
  CLKINVX1 U41 ( .A(A[53]), .Y(n15) );
  CLKINVX1 U42 ( .A(A[49]), .Y(n19) );
  CLKINVX1 U43 ( .A(A[41]), .Y(n27) );
  CLKINVX1 U44 ( .A(A[37]), .Y(n31) );
  CLKINVX1 U45 ( .A(A[33]), .Y(n35) );
  CLKINVX1 U46 ( .A(A[29]), .Y(n39) );
  CLKINVX1 U47 ( .A(A[25]), .Y(n43) );
  CLKINVX1 U48 ( .A(A[21]), .Y(n47) );
  CLKINVX1 U49 ( .A(A[17]), .Y(n51) );
  CLKINVX1 U50 ( .A(A[23]), .Y(n45) );
  CLKINVX1 U51 ( .A(A[19]), .Y(n49) );
  CLKINVX1 U52 ( .A(A[15]), .Y(n53) );
  CLKINVX1 U53 ( .A(A[11]), .Y(n57) );
  CLKINVX1 U54 ( .A(A[7]), .Y(n61) );
  CLKINVX1 U55 ( .A(A[3]), .Y(n65) );
  CLKINVX1 U56 ( .A(A[50]), .Y(n18) );
  CLKINVX1 U57 ( .A(A[24]), .Y(n44) );
  CLKINVX1 U58 ( .A(A[20]), .Y(n48) );
  CLKINVX1 U59 ( .A(A[16]), .Y(n52) );
  CLKINVX1 U60 ( .A(A[12]), .Y(n56) );
  CLKINVX1 U61 ( .A(A[8]), .Y(n60) );
  CLKINVX1 U62 ( .A(A[4]), .Y(n64) );
  CLKINVX1 U63 ( .A(A[10]), .Y(n58) );
  CLKINVX1 U64 ( .A(A[6]), .Y(n62) );
  CLKINVX1 U65 ( .A(A[13]), .Y(n55) );
  CLKINVX1 U66 ( .A(A[9]), .Y(n59) );
  CLKINVX1 U67 ( .A(A[5]), .Y(n63) );
  CLKINVX1 U68 ( .A(A[0]), .Y(n68) );
  CLKINVX1 U69 ( .A(A[1]), .Y(n67) );
  CLKMX2X2 U70 ( .A(A[9]), .B(AMUX1[9]), .S0(n3), .Y(ABSVAL[9]) );
  CLKMX2X2 U71 ( .A(A[8]), .B(AMUX1[8]), .S0(n4), .Y(ABSVAL[8]) );
  CLKMX2X2 U72 ( .A(A[7]), .B(AMUX1[7]), .S0(n4), .Y(ABSVAL[7]) );
  CLKMX2X2 U73 ( .A(A[6]), .B(AMUX1[6]), .S0(n4), .Y(ABSVAL[6]) );
  AND2X1 U74 ( .A(AMUX1[63]), .B(n4), .Y(ABSVAL[63]) );
  CLKMX2X2 U75 ( .A(A[62]), .B(AMUX1[62]), .S0(n4), .Y(ABSVAL[62]) );
  CLKMX2X2 U76 ( .A(A[60]), .B(AMUX1[60]), .S0(n4), .Y(ABSVAL[60]) );
  CLKMX2X2 U77 ( .A(A[5]), .B(AMUX1[5]), .S0(n4), .Y(ABSVAL[5]) );
  CLKMX2X2 U78 ( .A(A[59]), .B(AMUX1[59]), .S0(n4), .Y(ABSVAL[59]) );
  CLKMX2X2 U79 ( .A(A[58]), .B(AMUX1[58]), .S0(n4), .Y(ABSVAL[58]) );
  CLKMX2X2 U80 ( .A(A[57]), .B(AMUX1[57]), .S0(n4), .Y(ABSVAL[57]) );
  CLKMX2X2 U81 ( .A(A[56]), .B(AMUX1[56]), .S0(n3), .Y(ABSVAL[56]) );
  CLKMX2X2 U82 ( .A(A[55]), .B(AMUX1[55]), .S0(n3), .Y(ABSVAL[55]) );
  CLKMX2X2 U83 ( .A(A[54]), .B(AMUX1[54]), .S0(n3), .Y(ABSVAL[54]) );
  CLKMX2X2 U84 ( .A(A[53]), .B(AMUX1[53]), .S0(n3), .Y(ABSVAL[53]) );
  CLKMX2X2 U85 ( .A(A[52]), .B(AMUX1[52]), .S0(n3), .Y(ABSVAL[52]) );
  CLKMX2X2 U86 ( .A(A[51]), .B(AMUX1[51]), .S0(n3), .Y(ABSVAL[51]) );
  CLKMX2X2 U87 ( .A(A[50]), .B(AMUX1[50]), .S0(n3), .Y(ABSVAL[50]) );
  CLKMX2X2 U88 ( .A(A[4]), .B(AMUX1[4]), .S0(n3), .Y(ABSVAL[4]) );
  CLKMX2X2 U89 ( .A(A[49]), .B(AMUX1[49]), .S0(n3), .Y(ABSVAL[49]) );
  CLKMX2X2 U90 ( .A(A[48]), .B(AMUX1[48]), .S0(n3), .Y(ABSVAL[48]) );
  CLKMX2X2 U91 ( .A(A[47]), .B(AMUX1[47]), .S0(n3), .Y(ABSVAL[47]) );
  CLKMX2X2 U92 ( .A(A[46]), .B(AMUX1[46]), .S0(n3), .Y(ABSVAL[46]) );
  CLKMX2X2 U93 ( .A(A[45]), .B(AMUX1[45]), .S0(n3), .Y(ABSVAL[45]) );
  CLKMX2X2 U94 ( .A(A[44]), .B(AMUX1[44]), .S0(n2), .Y(ABSVAL[44]) );
  CLKMX2X2 U95 ( .A(A[43]), .B(AMUX1[43]), .S0(n2), .Y(ABSVAL[43]) );
  CLKMX2X2 U96 ( .A(A[42]), .B(AMUX1[42]), .S0(n2), .Y(ABSVAL[42]) );
  CLKMX2X2 U97 ( .A(A[41]), .B(AMUX1[41]), .S0(n2), .Y(ABSVAL[41]) );
  CLKMX2X2 U98 ( .A(A[40]), .B(AMUX1[40]), .S0(n2), .Y(ABSVAL[40]) );
  CLKMX2X2 U99 ( .A(A[3]), .B(AMUX1[3]), .S0(n2), .Y(ABSVAL[3]) );
  CLKMX2X2 U100 ( .A(A[39]), .B(AMUX1[39]), .S0(n2), .Y(ABSVAL[39]) );
  CLKMX2X2 U101 ( .A(A[38]), .B(AMUX1[38]), .S0(n2), .Y(ABSVAL[38]) );
  CLKMX2X2 U102 ( .A(A[37]), .B(AMUX1[37]), .S0(n2), .Y(ABSVAL[37]) );
  CLKMX2X2 U103 ( .A(A[36]), .B(AMUX1[36]), .S0(n2), .Y(ABSVAL[36]) );
  CLKMX2X2 U104 ( .A(A[35]), .B(AMUX1[35]), .S0(n2), .Y(ABSVAL[35]) );
  CLKMX2X2 U105 ( .A(A[34]), .B(AMUX1[34]), .S0(n2), .Y(ABSVAL[34]) );
  CLKMX2X2 U106 ( .A(A[33]), .B(AMUX1[33]), .S0(n1), .Y(ABSVAL[33]) );
  CLKMX2X2 U107 ( .A(A[32]), .B(AMUX1[32]), .S0(n1), .Y(ABSVAL[32]) );
  CLKMX2X2 U108 ( .A(A[31]), .B(AMUX1[31]), .S0(n1), .Y(ABSVAL[31]) );
  CLKMX2X2 U109 ( .A(A[30]), .B(AMUX1[30]), .S0(n1), .Y(ABSVAL[30]) );
  CLKMX2X2 U110 ( .A(A[2]), .B(AMUX1[2]), .S0(n1), .Y(ABSVAL[2]) );
  CLKMX2X2 U111 ( .A(A[29]), .B(AMUX1[29]), .S0(n1), .Y(ABSVAL[29]) );
  CLKMX2X2 U112 ( .A(A[28]), .B(AMUX1[28]), .S0(n1), .Y(ABSVAL[28]) );
  CLKMX2X2 U113 ( .A(A[27]), .B(AMUX1[27]), .S0(n1), .Y(ABSVAL[27]) );
  CLKMX2X2 U114 ( .A(A[26]), .B(AMUX1[26]), .S0(n1), .Y(ABSVAL[26]) );
  CLKMX2X2 U115 ( .A(A[25]), .B(AMUX1[25]), .S0(n1), .Y(ABSVAL[25]) );
  CLKMX2X2 U116 ( .A(A[24]), .B(AMUX1[24]), .S0(n1), .Y(ABSVAL[24]) );
  CLKMX2X2 U117 ( .A(A[23]), .B(AMUX1[23]), .S0(n1), .Y(ABSVAL[23]) );
  CLKMX2X2 U118 ( .A(A[22]), .B(AMUX1[22]), .S0(n1), .Y(ABSVAL[22]) );
  CLKMX2X2 U119 ( .A(A[21]), .B(AMUX1[21]), .S0(n1), .Y(ABSVAL[21]) );
  CLKMX2X2 U120 ( .A(A[20]), .B(AMUX1[20]), .S0(n1), .Y(ABSVAL[20]) );
  CLKMX2X2 U121 ( .A(A[19]), .B(AMUX1[19]), .S0(n1), .Y(ABSVAL[19]) );
  CLKMX2X2 U122 ( .A(A[18]), .B(AMUX1[18]), .S0(n1), .Y(ABSVAL[18]) );
  CLKMX2X2 U123 ( .A(A[17]), .B(AMUX1[17]), .S0(n2), .Y(ABSVAL[17]) );
  CLKMX2X2 U124 ( .A(A[16]), .B(AMUX1[16]), .S0(n2), .Y(ABSVAL[16]) );
  CLKMX2X2 U125 ( .A(A[15]), .B(AMUX1[15]), .S0(n2), .Y(ABSVAL[15]) );
  CLKMX2X2 U126 ( .A(A[14]), .B(AMUX1[14]), .S0(n2), .Y(ABSVAL[14]) );
  CLKMX2X2 U127 ( .A(A[13]), .B(AMUX1[13]), .S0(n3), .Y(ABSVAL[13]) );
  CLKMX2X2 U128 ( .A(A[12]), .B(AMUX1[12]), .S0(n3), .Y(ABSVAL[12]) );
  CLKMX2X2 U129 ( .A(A[11]), .B(AMUX1[11]), .S0(n3), .Y(ABSVAL[11]) );
  CLKMX2X2 U130 ( .A(A[10]), .B(AMUX1[10]), .S0(n2), .Y(ABSVAL[10]) );
endmodule


module GSIM_DW_inc_4 ( carry_in, a, carry_out, sum );
  input [63:0] a;
  output [63:0] sum;
  input carry_in;
  output carry_out;
  wire   \sum[63] , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63;
  assign sum[62] = \sum[63] ;
  assign sum[61] = \sum[63] ;
  assign sum[63] = \sum[63] ;

  ADDHXL U7 ( .A(a[59]), .B(n5), .CO(n4), .S(sum[59]) );
  ADDHXL U9 ( .A(a[57]), .B(n7), .CO(n6), .S(sum[57]) );
  ADDHXL U12 ( .A(a[54]), .B(n10), .CO(n9), .S(sum[54]) );
  ADDHXL U15 ( .A(a[51]), .B(n13), .CO(n12), .S(sum[51]) );
  ADDHXL U20 ( .A(a[46]), .B(n18), .CO(n17), .S(sum[46]) );
  ADDHXL U23 ( .A(a[43]), .B(n21), .CO(n20), .S(sum[43]) );
  ADDHXL U31 ( .A(a[35]), .B(n29), .CO(n28), .S(sum[35]) );
  ADDHXL U33 ( .A(a[33]), .B(n31), .CO(n30), .S(sum[33]) );
  ADDHXL U36 ( .A(a[30]), .B(n34), .CO(n33), .S(sum[30]) );
  ADDHXL U41 ( .A(a[25]), .B(n39), .CO(n38), .S(sum[25]) );
  ADDHXL U44 ( .A(a[22]), .B(n42), .CO(n41), .S(sum[22]) );
  ADDHXL U46 ( .A(a[20]), .B(n44), .CO(n43), .S(sum[20]) );
  ADDHXL U50 ( .A(a[16]), .B(n48), .CO(n47), .S(sum[16]) );
  ADDHXL U52 ( .A(a[14]), .B(n50), .CO(n49), .S(sum[14]) );
  ADDHXL U54 ( .A(a[12]), .B(n52), .CO(n51), .S(sum[12]) );
  ADDHXL U56 ( .A(a[10]), .B(n54), .CO(n53), .S(sum[10]) );
  ADDHXL U60 ( .A(a[6]), .B(n58), .CO(n57), .S(sum[6]) );
  ADDHXL U62 ( .A(a[4]), .B(n60), .CO(n59), .S(sum[4]) );
  ADDHXL U64 ( .A(a[2]), .B(n62), .CO(n61), .S(sum[2]) );
  ADDHXL U66 ( .A(carry_in), .B(a[0]), .CO(n63), .S(sum[0]) );
  ADDHXL U70 ( .A(a[11]), .B(n53), .CO(n52), .S(sum[11]) );
  ADDHXL U71 ( .A(a[13]), .B(n51), .CO(n50), .S(sum[13]) );
  ADDHXL U72 ( .A(a[15]), .B(n49), .CO(n48), .S(sum[15]) );
  ADDHXL U73 ( .A(a[17]), .B(n47), .CO(n46), .S(sum[17]) );
  ADDHXL U74 ( .A(a[19]), .B(n45), .CO(n44), .S(sum[19]) );
  ADDHXL U75 ( .A(a[23]), .B(n41), .CO(n40), .S(sum[23]) );
  ADDHXL U76 ( .A(a[21]), .B(n43), .CO(n42), .S(sum[21]) );
  ADDHXL U77 ( .A(a[1]), .B(n63), .CO(n62), .S(sum[1]) );
  ADDHXL U78 ( .A(a[5]), .B(n59), .CO(n58), .S(sum[5]) );
  ADDHXL U79 ( .A(a[9]), .B(n55), .CO(n54), .S(sum[9]) );
  ADDHXL U80 ( .A(a[3]), .B(n61), .CO(n60), .S(sum[3]) );
  ADDHXL U81 ( .A(a[7]), .B(n57), .CO(n56), .S(sum[7]) );
  ADDHXL U82 ( .A(a[26]), .B(n38), .CO(n37), .S(sum[26]) );
  ADDHXL U83 ( .A(a[29]), .B(n35), .CO(n34), .S(sum[29]) );
  ADDHXL U84 ( .A(a[31]), .B(n33), .CO(n32), .S(sum[31]) );
  ADDHXL U85 ( .A(a[34]), .B(n30), .CO(n29), .S(sum[34]) );
  ADDHXL U86 ( .A(a[36]), .B(n28), .CO(n27), .S(sum[36]) );
  ADDHXL U87 ( .A(a[39]), .B(n25), .CO(n24), .S(sum[39]) );
  ADDHXL U88 ( .A(a[41]), .B(n23), .CO(n22), .S(sum[41]) );
  ADDHXL U89 ( .A(a[44]), .B(n20), .CO(n19), .S(sum[44]) );
  ADDHXL U90 ( .A(a[47]), .B(n17), .CO(n16), .S(sum[47]) );
  ADDHXL U91 ( .A(a[48]), .B(n16), .CO(n15), .S(sum[48]) );
  ADDHXL U92 ( .A(a[50]), .B(n14), .CO(n13), .S(sum[50]) );
  ADDHXL U93 ( .A(a[52]), .B(n12), .CO(n11), .S(sum[52]) );
  ADDHXL U94 ( .A(a[55]), .B(n9), .CO(n8), .S(sum[55]) );
  ADDHXL U95 ( .A(a[56]), .B(n8), .CO(n7), .S(sum[56]) );
  ADDHXL U96 ( .A(a[58]), .B(n6), .CO(n5), .S(sum[58]) );
  ADDHXL U97 ( .A(a[53]), .B(n11), .CO(n10), .S(sum[53]) );
  ADDHXL U98 ( .A(a[42]), .B(n22), .CO(n21), .S(sum[42]) );
  ADDHXL U99 ( .A(a[24]), .B(n40), .CO(n39), .S(sum[24]) );
  ADDHXL U100 ( .A(a[37]), .B(n27), .CO(n26), .S(sum[37]) );
  ADDHXL U101 ( .A(a[40]), .B(n24), .CO(n23), .S(sum[40]) );
  ADDHXL U102 ( .A(a[32]), .B(n32), .CO(n31), .S(sum[32]) );
  ADDHXL U103 ( .A(a[27]), .B(n37), .CO(n36), .S(sum[27]) );
  ADDHXL U104 ( .A(a[45]), .B(n19), .CO(n18), .S(sum[45]) );
  NOR2BX1 U105 ( .AN(a[60]), .B(n4), .Y(\sum[63] ) );
  XOR2XL U106 ( .A(n4), .B(a[60]), .Y(sum[60]) );
  ADDHXL U107 ( .A(a[38]), .B(n26), .CO(n25), .S(sum[38]) );
  ADDHXL U108 ( .A(a[8]), .B(n56), .CO(n55), .S(sum[8]) );
  ADDHXL U109 ( .A(a[18]), .B(n46), .CO(n45), .S(sum[18]) );
  ADDHXL U110 ( .A(a[28]), .B(n36), .CO(n35), .S(sum[28]) );
  ADDHXL U111 ( .A(a[49]), .B(n15), .CO(n14), .S(sum[49]) );
endmodule


module GSIM_DW_div_tc_4 ( a, b, quotient, remainder, divide_by_0 );
  input [63:0] a;
  input [5:0] b;
  output [63:0] quotient;
  output [5:0] remainder;
  output divide_by_0;
  wire   \u_div/QInv[63] , \u_div/QInv[59] , \u_div/QInv[58] ,
         \u_div/QInv[57] , \u_div/QInv[56] , \u_div/QInv[55] ,
         \u_div/QInv[54] , \u_div/QInv[53] , \u_div/QInv[52] ,
         \u_div/QInv[51] , \u_div/QInv[50] , \u_div/QInv[49] ,
         \u_div/QInv[48] , \u_div/QInv[47] , \u_div/QInv[46] ,
         \u_div/QInv[45] , \u_div/QInv[44] , \u_div/QInv[43] ,
         \u_div/QInv[42] , \u_div/QInv[41] , \u_div/QInv[40] ,
         \u_div/QInv[39] , \u_div/QInv[38] , \u_div/QInv[37] ,
         \u_div/QInv[36] , \u_div/QInv[35] , \u_div/QInv[34] ,
         \u_div/QInv[33] , \u_div/QInv[32] , \u_div/QInv[31] ,
         \u_div/QInv[30] , \u_div/QInv[29] , \u_div/QInv[28] ,
         \u_div/QInv[27] , \u_div/QInv[26] , \u_div/QInv[25] ,
         \u_div/QInv[24] , \u_div/QInv[23] , \u_div/QInv[22] ,
         \u_div/QInv[21] , \u_div/QInv[20] , \u_div/QInv[19] ,
         \u_div/QInv[18] , \u_div/QInv[17] , \u_div/QInv[16] ,
         \u_div/QInv[15] , \u_div/QInv[14] , \u_div/QInv[13] ,
         \u_div/QInv[12] , \u_div/QInv[11] , \u_div/QInv[10] , \u_div/QInv[9] ,
         \u_div/QInv[8] , \u_div/QInv[7] , \u_div/QInv[6] , \u_div/QInv[5] ,
         \u_div/QInv[4] , \u_div/QInv[3] , \u_div/QInv[2] , \u_div/QInv[1] ,
         \u_div/QInv[0] , \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] ,
         \u_div/SumTmp[1][3] , \u_div/SumTmp[1][4] , \u_div/SumTmp[2][1] ,
         \u_div/SumTmp[2][2] , \u_div/SumTmp[2][3] , \u_div/SumTmp[2][4] ,
         \u_div/SumTmp[3][1] , \u_div/SumTmp[3][2] , \u_div/SumTmp[3][3] ,
         \u_div/SumTmp[3][4] , \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] ,
         \u_div/SumTmp[4][3] , \u_div/SumTmp[4][4] , \u_div/SumTmp[5][1] ,
         \u_div/SumTmp[5][2] , \u_div/SumTmp[5][3] , \u_div/SumTmp[5][4] ,
         \u_div/SumTmp[6][1] , \u_div/SumTmp[6][2] , \u_div/SumTmp[6][3] ,
         \u_div/SumTmp[6][4] , \u_div/SumTmp[7][1] , \u_div/SumTmp[7][2] ,
         \u_div/SumTmp[7][3] , \u_div/SumTmp[7][4] , \u_div/SumTmp[8][1] ,
         \u_div/SumTmp[8][2] , \u_div/SumTmp[8][3] , \u_div/SumTmp[8][4] ,
         \u_div/SumTmp[9][1] , \u_div/SumTmp[9][2] , \u_div/SumTmp[9][3] ,
         \u_div/SumTmp[9][4] , \u_div/SumTmp[10][1] , \u_div/SumTmp[10][2] ,
         \u_div/SumTmp[10][3] , \u_div/SumTmp[10][4] , \u_div/SumTmp[11][1] ,
         \u_div/SumTmp[11][2] , \u_div/SumTmp[11][3] , \u_div/SumTmp[11][4] ,
         \u_div/SumTmp[12][1] , \u_div/SumTmp[12][2] , \u_div/SumTmp[12][3] ,
         \u_div/SumTmp[12][4] , \u_div/SumTmp[13][1] , \u_div/SumTmp[13][2] ,
         \u_div/SumTmp[13][3] , \u_div/SumTmp[13][4] , \u_div/SumTmp[14][1] ,
         \u_div/SumTmp[14][2] , \u_div/SumTmp[14][3] , \u_div/SumTmp[14][4] ,
         \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] , \u_div/SumTmp[15][3] ,
         \u_div/SumTmp[15][4] , \u_div/SumTmp[16][1] , \u_div/SumTmp[16][2] ,
         \u_div/SumTmp[16][3] , \u_div/SumTmp[16][4] , \u_div/SumTmp[17][1] ,
         \u_div/SumTmp[17][2] , \u_div/SumTmp[17][3] , \u_div/SumTmp[17][4] ,
         \u_div/SumTmp[18][1] , \u_div/SumTmp[18][2] , \u_div/SumTmp[18][3] ,
         \u_div/SumTmp[18][4] , \u_div/SumTmp[19][1] , \u_div/SumTmp[19][2] ,
         \u_div/SumTmp[19][3] , \u_div/SumTmp[19][4] , \u_div/SumTmp[20][1] ,
         \u_div/SumTmp[20][2] , \u_div/SumTmp[20][3] , \u_div/SumTmp[20][4] ,
         \u_div/SumTmp[21][1] , \u_div/SumTmp[21][2] , \u_div/SumTmp[21][3] ,
         \u_div/SumTmp[21][4] , \u_div/SumTmp[22][1] , \u_div/SumTmp[22][2] ,
         \u_div/SumTmp[22][3] , \u_div/SumTmp[22][4] , \u_div/SumTmp[23][1] ,
         \u_div/SumTmp[23][2] , \u_div/SumTmp[23][3] , \u_div/SumTmp[23][4] ,
         \u_div/SumTmp[24][1] , \u_div/SumTmp[24][2] , \u_div/SumTmp[24][3] ,
         \u_div/SumTmp[24][4] , \u_div/SumTmp[25][1] , \u_div/SumTmp[25][2] ,
         \u_div/SumTmp[25][3] , \u_div/SumTmp[25][4] , \u_div/SumTmp[26][1] ,
         \u_div/SumTmp[26][2] , \u_div/SumTmp[26][3] , \u_div/SumTmp[26][4] ,
         \u_div/SumTmp[27][1] , \u_div/SumTmp[27][2] , \u_div/SumTmp[27][3] ,
         \u_div/SumTmp[27][4] , \u_div/SumTmp[28][1] , \u_div/SumTmp[28][2] ,
         \u_div/SumTmp[28][3] , \u_div/SumTmp[28][4] , \u_div/SumTmp[29][1] ,
         \u_div/SumTmp[29][2] , \u_div/SumTmp[29][3] , \u_div/SumTmp[29][4] ,
         \u_div/SumTmp[30][1] , \u_div/SumTmp[30][2] , \u_div/SumTmp[30][3] ,
         \u_div/SumTmp[30][4] , \u_div/SumTmp[31][1] , \u_div/SumTmp[31][2] ,
         \u_div/SumTmp[31][3] , \u_div/SumTmp[31][4] , \u_div/SumTmp[32][1] ,
         \u_div/SumTmp[32][2] , \u_div/SumTmp[32][3] , \u_div/SumTmp[32][4] ,
         \u_div/SumTmp[33][1] , \u_div/SumTmp[33][2] , \u_div/SumTmp[33][3] ,
         \u_div/SumTmp[33][4] , \u_div/SumTmp[34][1] , \u_div/SumTmp[34][2] ,
         \u_div/SumTmp[34][3] , \u_div/SumTmp[34][4] , \u_div/SumTmp[35][1] ,
         \u_div/SumTmp[35][2] , \u_div/SumTmp[35][3] , \u_div/SumTmp[35][4] ,
         \u_div/SumTmp[36][1] , \u_div/SumTmp[36][2] , \u_div/SumTmp[36][3] ,
         \u_div/SumTmp[36][4] , \u_div/SumTmp[37][1] , \u_div/SumTmp[37][2] ,
         \u_div/SumTmp[37][3] , \u_div/SumTmp[37][4] , \u_div/SumTmp[38][1] ,
         \u_div/SumTmp[38][2] , \u_div/SumTmp[38][3] , \u_div/SumTmp[38][4] ,
         \u_div/SumTmp[39][1] , \u_div/SumTmp[39][2] , \u_div/SumTmp[39][3] ,
         \u_div/SumTmp[39][4] , \u_div/SumTmp[40][1] , \u_div/SumTmp[40][2] ,
         \u_div/SumTmp[40][3] , \u_div/SumTmp[40][4] , \u_div/SumTmp[41][1] ,
         \u_div/SumTmp[41][2] , \u_div/SumTmp[41][3] , \u_div/SumTmp[41][4] ,
         \u_div/SumTmp[42][1] , \u_div/SumTmp[42][2] , \u_div/SumTmp[42][3] ,
         \u_div/SumTmp[42][4] , \u_div/SumTmp[43][1] , \u_div/SumTmp[43][2] ,
         \u_div/SumTmp[43][3] , \u_div/SumTmp[43][4] , \u_div/SumTmp[44][1] ,
         \u_div/SumTmp[44][2] , \u_div/SumTmp[44][3] , \u_div/SumTmp[44][4] ,
         \u_div/SumTmp[45][1] , \u_div/SumTmp[45][2] , \u_div/SumTmp[45][3] ,
         \u_div/SumTmp[45][4] , \u_div/SumTmp[46][1] , \u_div/SumTmp[46][2] ,
         \u_div/SumTmp[46][3] , \u_div/SumTmp[46][4] , \u_div/SumTmp[47][1] ,
         \u_div/SumTmp[47][2] , \u_div/SumTmp[47][3] , \u_div/SumTmp[47][4] ,
         \u_div/SumTmp[48][1] , \u_div/SumTmp[48][2] , \u_div/SumTmp[48][3] ,
         \u_div/SumTmp[48][4] , \u_div/SumTmp[49][1] , \u_div/SumTmp[49][2] ,
         \u_div/SumTmp[49][3] , \u_div/SumTmp[49][4] , \u_div/SumTmp[50][1] ,
         \u_div/SumTmp[50][2] , \u_div/SumTmp[50][3] , \u_div/SumTmp[50][4] ,
         \u_div/SumTmp[51][1] , \u_div/SumTmp[51][2] , \u_div/SumTmp[51][3] ,
         \u_div/SumTmp[51][4] , \u_div/SumTmp[52][1] , \u_div/SumTmp[52][2] ,
         \u_div/SumTmp[52][3] , \u_div/SumTmp[52][4] , \u_div/SumTmp[53][1] ,
         \u_div/SumTmp[53][2] , \u_div/SumTmp[53][3] , \u_div/SumTmp[53][4] ,
         \u_div/SumTmp[54][1] , \u_div/SumTmp[54][2] , \u_div/SumTmp[54][3] ,
         \u_div/SumTmp[54][4] , \u_div/SumTmp[55][1] , \u_div/SumTmp[55][2] ,
         \u_div/SumTmp[55][3] , \u_div/SumTmp[55][4] , \u_div/SumTmp[56][1] ,
         \u_div/SumTmp[56][2] , \u_div/SumTmp[56][3] , \u_div/SumTmp[56][4] ,
         \u_div/SumTmp[57][1] , \u_div/SumTmp[57][2] , \u_div/SumTmp[57][3] ,
         \u_div/SumTmp[57][4] , \u_div/SumTmp[58][1] , \u_div/SumTmp[58][2] ,
         \u_div/SumTmp[58][3] , \u_div/SumTmp[58][4] , \u_div/SumTmp[59][3] ,
         \u_div/SumTmp[59][4] , \u_div/CryTmp[0][6] , \u_div/CryTmp[1][6] ,
         \u_div/CryTmp[2][6] , \u_div/CryTmp[3][6] , \u_div/CryTmp[4][6] ,
         \u_div/CryTmp[5][6] , \u_div/CryTmp[6][6] , \u_div/CryTmp[7][6] ,
         \u_div/CryTmp[8][6] , \u_div/CryTmp[9][6] , \u_div/CryTmp[10][6] ,
         \u_div/CryTmp[11][6] , \u_div/CryTmp[12][6] , \u_div/CryTmp[13][6] ,
         \u_div/CryTmp[14][6] , \u_div/CryTmp[15][6] , \u_div/CryTmp[16][6] ,
         \u_div/CryTmp[17][6] , \u_div/CryTmp[18][6] , \u_div/CryTmp[19][6] ,
         \u_div/CryTmp[20][6] , \u_div/CryTmp[21][6] , \u_div/CryTmp[22][6] ,
         \u_div/CryTmp[23][6] , \u_div/CryTmp[24][6] , \u_div/CryTmp[25][6] ,
         \u_div/CryTmp[26][6] , \u_div/CryTmp[27][6] , \u_div/CryTmp[28][6] ,
         \u_div/CryTmp[29][6] , \u_div/CryTmp[30][6] , \u_div/CryTmp[31][6] ,
         \u_div/CryTmp[32][6] , \u_div/CryTmp[33][6] , \u_div/CryTmp[34][6] ,
         \u_div/CryTmp[35][6] , \u_div/CryTmp[36][6] , \u_div/CryTmp[37][6] ,
         \u_div/CryTmp[38][6] , \u_div/CryTmp[39][6] , \u_div/CryTmp[40][6] ,
         \u_div/CryTmp[41][6] , \u_div/CryTmp[42][6] , \u_div/CryTmp[43][6] ,
         \u_div/CryTmp[44][6] , \u_div/CryTmp[45][6] , \u_div/CryTmp[46][6] ,
         \u_div/CryTmp[47][6] , \u_div/CryTmp[48][6] , \u_div/CryTmp[49][6] ,
         \u_div/CryTmp[50][6] , \u_div/CryTmp[51][6] , \u_div/CryTmp[52][6] ,
         \u_div/CryTmp[53][6] , \u_div/CryTmp[54][6] , \u_div/CryTmp[55][6] ,
         \u_div/CryTmp[56][6] , \u_div/CryTmp[57][6] , \u_div/CryTmp[58][6] ,
         \u_div/CryTmp[59][6] , \u_div/PartRem[1][3] , \u_div/PartRem[1][4] ,
         \u_div/PartRem[1][5] , \u_div/PartRem[2][2] , \u_div/PartRem[2][3] ,
         \u_div/PartRem[2][4] , \u_div/PartRem[2][5] , \u_div/PartRem[3][0] ,
         \u_div/PartRem[3][2] , \u_div/PartRem[3][3] , \u_div/PartRem[3][4] ,
         \u_div/PartRem[3][5] , \u_div/PartRem[4][0] , \u_div/PartRem[4][2] ,
         \u_div/PartRem[4][3] , \u_div/PartRem[4][4] , \u_div/PartRem[4][5] ,
         \u_div/PartRem[5][0] , \u_div/PartRem[5][2] , \u_div/PartRem[5][3] ,
         \u_div/PartRem[5][4] , \u_div/PartRem[5][5] , \u_div/PartRem[6][0] ,
         \u_div/PartRem[6][2] , \u_div/PartRem[6][3] , \u_div/PartRem[6][4] ,
         \u_div/PartRem[6][5] , \u_div/PartRem[7][0] , \u_div/PartRem[7][2] ,
         \u_div/PartRem[7][3] , \u_div/PartRem[7][4] , \u_div/PartRem[7][5] ,
         \u_div/PartRem[8][0] , \u_div/PartRem[8][2] , \u_div/PartRem[8][3] ,
         \u_div/PartRem[8][4] , \u_div/PartRem[8][5] , \u_div/PartRem[9][0] ,
         \u_div/PartRem[9][2] , \u_div/PartRem[9][3] , \u_div/PartRem[9][4] ,
         \u_div/PartRem[9][5] , \u_div/PartRem[10][0] , \u_div/PartRem[10][2] ,
         \u_div/PartRem[10][3] , \u_div/PartRem[10][4] ,
         \u_div/PartRem[10][5] , \u_div/PartRem[11][0] ,
         \u_div/PartRem[11][2] , \u_div/PartRem[11][3] ,
         \u_div/PartRem[11][4] , \u_div/PartRem[11][5] ,
         \u_div/PartRem[12][0] , \u_div/PartRem[12][2] ,
         \u_div/PartRem[12][3] , \u_div/PartRem[12][4] ,
         \u_div/PartRem[12][5] , \u_div/PartRem[13][0] ,
         \u_div/PartRem[13][2] , \u_div/PartRem[13][3] ,
         \u_div/PartRem[13][4] , \u_div/PartRem[13][5] ,
         \u_div/PartRem[14][0] , \u_div/PartRem[14][2] ,
         \u_div/PartRem[14][3] , \u_div/PartRem[14][4] ,
         \u_div/PartRem[14][5] , \u_div/PartRem[15][0] ,
         \u_div/PartRem[15][2] , \u_div/PartRem[15][3] ,
         \u_div/PartRem[15][4] , \u_div/PartRem[15][5] ,
         \u_div/PartRem[16][0] , \u_div/PartRem[16][2] ,
         \u_div/PartRem[16][3] , \u_div/PartRem[16][4] ,
         \u_div/PartRem[16][5] , \u_div/PartRem[17][0] ,
         \u_div/PartRem[17][2] , \u_div/PartRem[17][3] ,
         \u_div/PartRem[17][4] , \u_div/PartRem[17][5] ,
         \u_div/PartRem[18][0] , \u_div/PartRem[18][2] ,
         \u_div/PartRem[18][3] , \u_div/PartRem[18][4] ,
         \u_div/PartRem[18][5] , \u_div/PartRem[19][0] ,
         \u_div/PartRem[19][2] , \u_div/PartRem[19][3] ,
         \u_div/PartRem[19][4] , \u_div/PartRem[19][5] ,
         \u_div/PartRem[20][0] , \u_div/PartRem[20][2] ,
         \u_div/PartRem[20][3] , \u_div/PartRem[20][4] ,
         \u_div/PartRem[20][5] , \u_div/PartRem[21][0] ,
         \u_div/PartRem[21][2] , \u_div/PartRem[21][3] ,
         \u_div/PartRem[21][4] , \u_div/PartRem[21][5] ,
         \u_div/PartRem[22][0] , \u_div/PartRem[22][2] ,
         \u_div/PartRem[22][3] , \u_div/PartRem[22][4] ,
         \u_div/PartRem[22][5] , \u_div/PartRem[23][0] ,
         \u_div/PartRem[23][2] , \u_div/PartRem[23][3] ,
         \u_div/PartRem[23][4] , \u_div/PartRem[23][5] ,
         \u_div/PartRem[24][0] , \u_div/PartRem[24][2] ,
         \u_div/PartRem[24][3] , \u_div/PartRem[24][4] ,
         \u_div/PartRem[24][5] , \u_div/PartRem[25][0] ,
         \u_div/PartRem[25][2] , \u_div/PartRem[25][3] ,
         \u_div/PartRem[25][4] , \u_div/PartRem[25][5] ,
         \u_div/PartRem[26][0] , \u_div/PartRem[26][2] ,
         \u_div/PartRem[26][3] , \u_div/PartRem[26][4] ,
         \u_div/PartRem[26][5] , \u_div/PartRem[27][0] ,
         \u_div/PartRem[27][2] , \u_div/PartRem[27][3] ,
         \u_div/PartRem[27][4] , \u_div/PartRem[27][5] ,
         \u_div/PartRem[28][0] , \u_div/PartRem[28][2] ,
         \u_div/PartRem[28][3] , \u_div/PartRem[28][4] ,
         \u_div/PartRem[28][5] , \u_div/PartRem[29][0] ,
         \u_div/PartRem[29][2] , \u_div/PartRem[29][3] ,
         \u_div/PartRem[29][4] , \u_div/PartRem[29][5] ,
         \u_div/PartRem[30][0] , \u_div/PartRem[30][2] ,
         \u_div/PartRem[30][3] , \u_div/PartRem[30][4] ,
         \u_div/PartRem[30][5] , \u_div/PartRem[31][0] ,
         \u_div/PartRem[31][2] , \u_div/PartRem[31][3] ,
         \u_div/PartRem[31][4] , \u_div/PartRem[31][5] ,
         \u_div/PartRem[32][0] , \u_div/PartRem[32][2] ,
         \u_div/PartRem[32][3] , \u_div/PartRem[32][4] ,
         \u_div/PartRem[32][5] , \u_div/PartRem[33][0] ,
         \u_div/PartRem[33][2] , \u_div/PartRem[33][3] ,
         \u_div/PartRem[33][4] , \u_div/PartRem[33][5] ,
         \u_div/PartRem[34][0] , \u_div/PartRem[34][2] ,
         \u_div/PartRem[34][3] , \u_div/PartRem[34][4] ,
         \u_div/PartRem[34][5] , \u_div/PartRem[35][0] ,
         \u_div/PartRem[35][2] , \u_div/PartRem[35][3] ,
         \u_div/PartRem[35][4] , \u_div/PartRem[35][5] ,
         \u_div/PartRem[36][0] , \u_div/PartRem[36][2] ,
         \u_div/PartRem[36][3] , \u_div/PartRem[36][4] ,
         \u_div/PartRem[36][5] , \u_div/PartRem[37][0] ,
         \u_div/PartRem[37][2] , \u_div/PartRem[37][3] ,
         \u_div/PartRem[37][4] , \u_div/PartRem[37][5] ,
         \u_div/PartRem[38][0] , \u_div/PartRem[38][2] ,
         \u_div/PartRem[38][3] , \u_div/PartRem[38][4] ,
         \u_div/PartRem[38][5] , \u_div/PartRem[39][0] ,
         \u_div/PartRem[39][2] , \u_div/PartRem[39][3] ,
         \u_div/PartRem[39][4] , \u_div/PartRem[39][5] ,
         \u_div/PartRem[40][0] , \u_div/PartRem[40][2] ,
         \u_div/PartRem[40][3] , \u_div/PartRem[40][4] ,
         \u_div/PartRem[40][5] , \u_div/PartRem[41][0] ,
         \u_div/PartRem[41][2] , \u_div/PartRem[41][3] ,
         \u_div/PartRem[41][4] , \u_div/PartRem[41][5] ,
         \u_div/PartRem[42][0] , \u_div/PartRem[42][2] ,
         \u_div/PartRem[42][3] , \u_div/PartRem[42][4] ,
         \u_div/PartRem[42][5] , \u_div/PartRem[43][0] ,
         \u_div/PartRem[43][2] , \u_div/PartRem[43][3] ,
         \u_div/PartRem[43][4] , \u_div/PartRem[43][5] ,
         \u_div/PartRem[44][0] , \u_div/PartRem[44][2] ,
         \u_div/PartRem[44][3] , \u_div/PartRem[44][4] ,
         \u_div/PartRem[44][5] , \u_div/PartRem[45][0] ,
         \u_div/PartRem[45][2] , \u_div/PartRem[45][3] ,
         \u_div/PartRem[45][4] , \u_div/PartRem[45][5] ,
         \u_div/PartRem[46][0] , \u_div/PartRem[46][2] ,
         \u_div/PartRem[46][3] , \u_div/PartRem[46][4] ,
         \u_div/PartRem[46][5] , \u_div/PartRem[47][0] ,
         \u_div/PartRem[47][2] , \u_div/PartRem[47][3] ,
         \u_div/PartRem[47][4] , \u_div/PartRem[47][5] ,
         \u_div/PartRem[48][0] , \u_div/PartRem[48][2] ,
         \u_div/PartRem[48][3] , \u_div/PartRem[48][4] ,
         \u_div/PartRem[48][5] , \u_div/PartRem[49][0] ,
         \u_div/PartRem[49][2] , \u_div/PartRem[49][3] ,
         \u_div/PartRem[49][4] , \u_div/PartRem[49][5] ,
         \u_div/PartRem[50][0] , \u_div/PartRem[50][2] ,
         \u_div/PartRem[50][3] , \u_div/PartRem[50][4] ,
         \u_div/PartRem[50][5] , \u_div/PartRem[51][0] ,
         \u_div/PartRem[51][2] , \u_div/PartRem[51][3] ,
         \u_div/PartRem[51][4] , \u_div/PartRem[51][5] ,
         \u_div/PartRem[52][0] , \u_div/PartRem[52][2] ,
         \u_div/PartRem[52][3] , \u_div/PartRem[52][4] ,
         \u_div/PartRem[52][5] , \u_div/PartRem[53][0] ,
         \u_div/PartRem[53][2] , \u_div/PartRem[53][3] ,
         \u_div/PartRem[53][4] , \u_div/PartRem[53][5] ,
         \u_div/PartRem[54][0] , \u_div/PartRem[54][2] ,
         \u_div/PartRem[54][3] , \u_div/PartRem[54][4] ,
         \u_div/PartRem[54][5] , \u_div/PartRem[55][0] ,
         \u_div/PartRem[55][2] , \u_div/PartRem[55][3] ,
         \u_div/PartRem[55][4] , \u_div/PartRem[55][5] ,
         \u_div/PartRem[56][0] , \u_div/PartRem[56][2] ,
         \u_div/PartRem[56][3] , \u_div/PartRem[56][4] ,
         \u_div/PartRem[56][5] , \u_div/PartRem[57][0] ,
         \u_div/PartRem[57][2] , \u_div/PartRem[57][3] ,
         \u_div/PartRem[57][4] , \u_div/PartRem[57][5] ,
         \u_div/PartRem[58][0] , \u_div/PartRem[58][2] ,
         \u_div/PartRem[58][3] , \u_div/PartRem[58][4] ,
         \u_div/PartRem[58][5] , \u_div/PartRem[59][0] ,
         \u_div/PartRem[59][2] , \u_div/PartRem[59][3] ,
         \u_div/PartRem[59][4] , \u_div/PartRem[59][5] ,
         \u_div/PartRem[60][0] , \u_div/PartRem[61][0] ,
         \u_div/PartRem[62][0] , \u_div/PartRem[63][0] ,
         \u_div/PartRem[64][0] , \u_div/u_add_PartRem_2_1/n3 ,
         \u_div/u_add_PartRem_2_1/n2 , \u_div/u_add_PartRem_2_2/n3 ,
         \u_div/u_add_PartRem_2_2/n2 , \u_div/u_add_PartRem_2_3/n3 ,
         \u_div/u_add_PartRem_2_3/n2 , \u_div/u_add_PartRem_2_4/n3 ,
         \u_div/u_add_PartRem_2_4/n2 , \u_div/u_add_PartRem_2_5/n3 ,
         \u_div/u_add_PartRem_2_5/n2 , \u_div/u_add_PartRem_2_6/n3 ,
         \u_div/u_add_PartRem_2_6/n2 , \u_div/u_add_PartRem_2_7/n3 ,
         \u_div/u_add_PartRem_2_7/n2 , \u_div/u_add_PartRem_2_8/n3 ,
         \u_div/u_add_PartRem_2_8/n2 , \u_div/u_add_PartRem_2_9/n3 ,
         \u_div/u_add_PartRem_2_9/n2 , \u_div/u_add_PartRem_2_10/n3 ,
         \u_div/u_add_PartRem_2_10/n2 , \u_div/u_add_PartRem_2_11/n3 ,
         \u_div/u_add_PartRem_2_11/n2 , \u_div/u_add_PartRem_2_12/n3 ,
         \u_div/u_add_PartRem_2_12/n2 , \u_div/u_add_PartRem_2_13/n3 ,
         \u_div/u_add_PartRem_2_13/n2 , \u_div/u_add_PartRem_2_14/n3 ,
         \u_div/u_add_PartRem_2_14/n2 , \u_div/u_add_PartRem_2_15/n3 ,
         \u_div/u_add_PartRem_2_15/n2 , \u_div/u_add_PartRem_2_16/n3 ,
         \u_div/u_add_PartRem_2_16/n2 , \u_div/u_add_PartRem_2_17/n3 ,
         \u_div/u_add_PartRem_2_17/n2 , \u_div/u_add_PartRem_2_18/n3 ,
         \u_div/u_add_PartRem_2_18/n2 , \u_div/u_add_PartRem_2_19/n3 ,
         \u_div/u_add_PartRem_2_19/n2 , \u_div/u_add_PartRem_2_20/n3 ,
         \u_div/u_add_PartRem_2_20/n2 , \u_div/u_add_PartRem_2_21/n3 ,
         \u_div/u_add_PartRem_2_21/n2 , \u_div/u_add_PartRem_2_22/n3 ,
         \u_div/u_add_PartRem_2_22/n2 , \u_div/u_add_PartRem_2_23/n3 ,
         \u_div/u_add_PartRem_2_23/n2 , \u_div/u_add_PartRem_2_24/n3 ,
         \u_div/u_add_PartRem_2_24/n2 , \u_div/u_add_PartRem_2_25/n3 ,
         \u_div/u_add_PartRem_2_25/n2 , \u_div/u_add_PartRem_2_26/n3 ,
         \u_div/u_add_PartRem_2_26/n2 , \u_div/u_add_PartRem_2_27/n3 ,
         \u_div/u_add_PartRem_2_27/n2 , \u_div/u_add_PartRem_2_28/n3 ,
         \u_div/u_add_PartRem_2_28/n2 , \u_div/u_add_PartRem_2_29/n3 ,
         \u_div/u_add_PartRem_2_29/n2 , \u_div/u_add_PartRem_2_30/n3 ,
         \u_div/u_add_PartRem_2_30/n2 , \u_div/u_add_PartRem_2_31/n3 ,
         \u_div/u_add_PartRem_2_31/n2 , \u_div/u_add_PartRem_2_32/n3 ,
         \u_div/u_add_PartRem_2_32/n2 , \u_div/u_add_PartRem_2_33/n3 ,
         \u_div/u_add_PartRem_2_33/n2 , \u_div/u_add_PartRem_2_34/n3 ,
         \u_div/u_add_PartRem_2_34/n2 , \u_div/u_add_PartRem_2_35/n3 ,
         \u_div/u_add_PartRem_2_35/n2 , \u_div/u_add_PartRem_2_36/n3 ,
         \u_div/u_add_PartRem_2_36/n2 , \u_div/u_add_PartRem_2_37/n3 ,
         \u_div/u_add_PartRem_2_37/n2 , \u_div/u_add_PartRem_2_38/n3 ,
         \u_div/u_add_PartRem_2_38/n2 , \u_div/u_add_PartRem_2_39/n3 ,
         \u_div/u_add_PartRem_2_39/n2 , \u_div/u_add_PartRem_2_40/n3 ,
         \u_div/u_add_PartRem_2_40/n2 , \u_div/u_add_PartRem_2_41/n3 ,
         \u_div/u_add_PartRem_2_41/n2 , \u_div/u_add_PartRem_2_42/n3 ,
         \u_div/u_add_PartRem_2_42/n2 , \u_div/u_add_PartRem_2_43/n3 ,
         \u_div/u_add_PartRem_2_43/n2 , \u_div/u_add_PartRem_2_44/n3 ,
         \u_div/u_add_PartRem_2_44/n2 , \u_div/u_add_PartRem_2_45/n3 ,
         \u_div/u_add_PartRem_2_45/n2 , \u_div/u_add_PartRem_2_46/n3 ,
         \u_div/u_add_PartRem_2_46/n2 , \u_div/u_add_PartRem_2_47/n3 ,
         \u_div/u_add_PartRem_2_47/n2 , \u_div/u_add_PartRem_2_48/n3 ,
         \u_div/u_add_PartRem_2_48/n2 , \u_div/u_add_PartRem_2_49/n3 ,
         \u_div/u_add_PartRem_2_49/n2 , \u_div/u_add_PartRem_2_50/n3 ,
         \u_div/u_add_PartRem_2_50/n2 , \u_div/u_add_PartRem_2_51/n3 ,
         \u_div/u_add_PartRem_2_51/n2 , \u_div/u_add_PartRem_2_52/n3 ,
         \u_div/u_add_PartRem_2_52/n2 , \u_div/u_add_PartRem_2_53/n3 ,
         \u_div/u_add_PartRem_2_53/n2 , \u_div/u_add_PartRem_2_54/n3 ,
         \u_div/u_add_PartRem_2_54/n2 , \u_div/u_add_PartRem_2_55/n3 ,
         \u_div/u_add_PartRem_2_55/n2 , \u_div/u_add_PartRem_2_56/n3 ,
         \u_div/u_add_PartRem_2_56/n2 , \u_div/u_add_PartRem_2_57/n3 ,
         \u_div/u_add_PartRem_2_57/n2 , \u_div/u_add_PartRem_2_58/n3 ,
         \u_div/u_add_PartRem_2_58/n2 , n1, n2, n3, n4, n5, n6, n7, n8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign \u_div/QInv[63]  = a[63];

  GSIM_DW01_absval_4 \u_div/u_absval_AAbs  ( .A({n3, a[62:0]}), .ABSVAL({
        \u_div/PartRem[64][0] , \u_div/PartRem[63][0] , \u_div/PartRem[62][0] , 
        \u_div/PartRem[61][0] , \u_div/PartRem[60][0] , \u_div/PartRem[59][0] , 
        \u_div/PartRem[58][0] , \u_div/PartRem[57][0] , \u_div/PartRem[56][0] , 
        \u_div/PartRem[55][0] , \u_div/PartRem[54][0] , \u_div/PartRem[53][0] , 
        \u_div/PartRem[52][0] , \u_div/PartRem[51][0] , \u_div/PartRem[50][0] , 
        \u_div/PartRem[49][0] , \u_div/PartRem[48][0] , \u_div/PartRem[47][0] , 
        \u_div/PartRem[46][0] , \u_div/PartRem[45][0] , \u_div/PartRem[44][0] , 
        \u_div/PartRem[43][0] , \u_div/PartRem[42][0] , \u_div/PartRem[41][0] , 
        \u_div/PartRem[40][0] , \u_div/PartRem[39][0] , \u_div/PartRem[38][0] , 
        \u_div/PartRem[37][0] , \u_div/PartRem[36][0] , \u_div/PartRem[35][0] , 
        \u_div/PartRem[34][0] , \u_div/PartRem[33][0] , \u_div/PartRem[32][0] , 
        \u_div/PartRem[31][0] , \u_div/PartRem[30][0] , \u_div/PartRem[29][0] , 
        \u_div/PartRem[28][0] , \u_div/PartRem[27][0] , \u_div/PartRem[26][0] , 
        \u_div/PartRem[25][0] , \u_div/PartRem[24][0] , \u_div/PartRem[23][0] , 
        \u_div/PartRem[22][0] , \u_div/PartRem[21][0] , \u_div/PartRem[20][0] , 
        \u_div/PartRem[19][0] , \u_div/PartRem[18][0] , \u_div/PartRem[17][0] , 
        \u_div/PartRem[16][0] , \u_div/PartRem[15][0] , \u_div/PartRem[14][0] , 
        \u_div/PartRem[13][0] , \u_div/PartRem[12][0] , \u_div/PartRem[11][0] , 
        \u_div/PartRem[10][0] , \u_div/PartRem[9][0] , \u_div/PartRem[8][0] , 
        \u_div/PartRem[7][0] , \u_div/PartRem[6][0] , \u_div/PartRem[5][0] , 
        \u_div/PartRem[4][0] , \u_div/PartRem[3][0] , SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1}) );
  GSIM_DW_inc_4 \u_div/u_inc_QInc  ( .carry_in(n4), .a({n3, n3, n3, 
        \u_div/QInv[63] , \u_div/QInv[59] , \u_div/QInv[58] , \u_div/QInv[57] , 
        \u_div/QInv[56] , \u_div/QInv[55] , \u_div/QInv[54] , \u_div/QInv[53] , 
        \u_div/QInv[52] , \u_div/QInv[51] , \u_div/QInv[50] , \u_div/QInv[49] , 
        \u_div/QInv[48] , \u_div/QInv[47] , \u_div/QInv[46] , \u_div/QInv[45] , 
        \u_div/QInv[44] , \u_div/QInv[43] , \u_div/QInv[42] , \u_div/QInv[41] , 
        \u_div/QInv[40] , \u_div/QInv[39] , \u_div/QInv[38] , \u_div/QInv[37] , 
        \u_div/QInv[36] , \u_div/QInv[35] , \u_div/QInv[34] , \u_div/QInv[33] , 
        \u_div/QInv[32] , \u_div/QInv[31] , \u_div/QInv[30] , \u_div/QInv[29] , 
        \u_div/QInv[28] , \u_div/QInv[27] , \u_div/QInv[26] , \u_div/QInv[25] , 
        \u_div/QInv[24] , \u_div/QInv[23] , \u_div/QInv[22] , \u_div/QInv[21] , 
        \u_div/QInv[20] , \u_div/QInv[19] , \u_div/QInv[18] , \u_div/QInv[17] , 
        \u_div/QInv[16] , \u_div/QInv[15] , \u_div/QInv[14] , \u_div/QInv[13] , 
        \u_div/QInv[12] , \u_div/QInv[11] , \u_div/QInv[10] , \u_div/QInv[9] , 
        \u_div/QInv[8] , \u_div/QInv[7] , \u_div/QInv[6] , \u_div/QInv[5] , 
        \u_div/QInv[4] , \u_div/QInv[3] , \u_div/QInv[2] , \u_div/QInv[1] , 
        \u_div/QInv[0] }), .sum(quotient) );
  MX2XL \u_div/u_mx_PartRem_1_2_0  ( .A(\u_div/PartRem[3][0] ), .B(
        \u_div/PartRem[3][0] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/SumTmp[1][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_0  ( .A(\u_div/PartRem[7][0] ), .B(
        \u_div/PartRem[7][0] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/SumTmp[5][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_5_1  ( .A(\u_div/SumTmp[5][1] ), .B(
        \u_div/SumTmp[5][1] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_0  ( .A(\u_div/PartRem[12][0] ), .B(
        \u_div/PartRem[12][0] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/SumTmp[10][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_10_1  ( .A(\u_div/SumTmp[10][1] ), .B(
        \u_div/SumTmp[10][1] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_0  ( .A(\u_div/PartRem[17][0] ), .B(
        \u_div/PartRem[17][0] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/SumTmp[15][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_15_1  ( .A(\u_div/SumTmp[15][1] ), .B(
        \u_div/SumTmp[15][1] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_0  ( .A(\u_div/PartRem[22][0] ), .B(
        \u_div/PartRem[22][0] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/SumTmp[20][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_20_1  ( .A(\u_div/SumTmp[20][1] ), .B(
        \u_div/SumTmp[20][1] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_0  ( .A(\u_div/PartRem[27][0] ), .B(
        \u_div/PartRem[27][0] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/SumTmp[25][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_25_1  ( .A(\u_div/SumTmp[25][1] ), .B(
        \u_div/SumTmp[25][1] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_0  ( .A(\u_div/PartRem[32][0] ), .B(
        \u_div/PartRem[32][0] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/SumTmp[30][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_30_1  ( .A(\u_div/SumTmp[30][1] ), .B(
        \u_div/SumTmp[30][1] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_0  ( .A(\u_div/PartRem[37][0] ), .B(
        \u_div/PartRem[37][0] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/SumTmp[35][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_35_1  ( .A(\u_div/SumTmp[35][1] ), .B(
        \u_div/SumTmp[35][1] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_0  ( .A(\u_div/PartRem[42][0] ), .B(
        \u_div/PartRem[42][0] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/SumTmp[40][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_40_1  ( .A(\u_div/SumTmp[40][1] ), .B(
        \u_div/SumTmp[40][1] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_0  ( .A(\u_div/PartRem[47][0] ), .B(
        \u_div/PartRem[47][0] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/SumTmp[45][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_45_1  ( .A(\u_div/SumTmp[45][1] ), .B(
        \u_div/SumTmp[45][1] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_0  ( .A(\u_div/PartRem[52][0] ), .B(
        \u_div/PartRem[52][0] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/SumTmp[50][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_50_1  ( .A(\u_div/SumTmp[50][1] ), .B(
        \u_div/SumTmp[50][1] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_55_1  ( .A(\u_div/SumTmp[55][1] ), .B(
        \u_div/SumTmp[55][1] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_0  ( .A(\u_div/PartRem[4][0] ), .B(
        \u_div/PartRem[4][0] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/SumTmp[2][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_0  ( .A(\u_div/PartRem[5][0] ), .B(
        \u_div/PartRem[5][0] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/SumTmp[3][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_0  ( .A(\u_div/PartRem[8][0] ), .B(
        \u_div/PartRem[8][0] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/SumTmp[6][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_0  ( .A(\u_div/PartRem[13][0] ), .B(
        \u_div/PartRem[13][0] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/SumTmp[11][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_0  ( .A(\u_div/PartRem[14][0] ), .B(
        \u_div/PartRem[14][0] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/SumTmp[12][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_0  ( .A(\u_div/PartRem[15][0] ), .B(
        \u_div/PartRem[15][0] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/SumTmp[13][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_0  ( .A(\u_div/PartRem[18][0] ), .B(
        \u_div/PartRem[18][0] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/SumTmp[16][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_0  ( .A(\u_div/PartRem[19][0] ), .B(
        \u_div/PartRem[19][0] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/SumTmp[17][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_0  ( .A(\u_div/PartRem[23][0] ), .B(
        \u_div/PartRem[23][0] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/SumTmp[21][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_0  ( .A(\u_div/PartRem[24][0] ), .B(
        \u_div/PartRem[24][0] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/SumTmp[22][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_0  ( .A(\u_div/PartRem[25][0] ), .B(
        \u_div/PartRem[25][0] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/SumTmp[23][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_0  ( .A(\u_div/PartRem[28][0] ), .B(
        \u_div/PartRem[28][0] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/SumTmp[26][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_0  ( .A(\u_div/PartRem[30][0] ), .B(
        \u_div/PartRem[30][0] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/SumTmp[28][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_0  ( .A(\u_div/PartRem[33][0] ), .B(
        \u_div/PartRem[33][0] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/SumTmp[31][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_0  ( .A(\u_div/PartRem[34][0] ), .B(
        \u_div/PartRem[34][0] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/SumTmp[32][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_0  ( .A(\u_div/PartRem[35][0] ), .B(
        \u_div/PartRem[35][0] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/SumTmp[33][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_0  ( .A(\u_div/PartRem[38][0] ), .B(
        \u_div/PartRem[38][0] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/SumTmp[36][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_0  ( .A(\u_div/PartRem[40][0] ), .B(
        \u_div/PartRem[40][0] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/SumTmp[38][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_0  ( .A(\u_div/PartRem[43][0] ), .B(
        \u_div/PartRem[43][0] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/SumTmp[41][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_0  ( .A(\u_div/PartRem[44][0] ), .B(
        \u_div/PartRem[44][0] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/SumTmp[42][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_0  ( .A(\u_div/PartRem[45][0] ), .B(
        \u_div/PartRem[45][0] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/SumTmp[43][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_0  ( .A(\u_div/PartRem[48][0] ), .B(
        \u_div/PartRem[48][0] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/SumTmp[46][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_0  ( .A(\u_div/PartRem[53][0] ), .B(
        \u_div/PartRem[53][0] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/SumTmp[51][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_0  ( .A(\u_div/PartRem[54][0] ), .B(
        \u_div/PartRem[54][0] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/SumTmp[52][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_0  ( .A(\u_div/PartRem[55][0] ), .B(
        \u_div/PartRem[55][0] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/SumTmp[53][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_0  ( .A(\u_div/PartRem[58][0] ), .B(
        \u_div/PartRem[58][0] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/SumTmp[56][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_0  ( .A(\u_div/PartRem[59][0] ), .B(
        \u_div/PartRem[59][0] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/SumTmp[57][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_0  ( .A(\u_div/PartRem[60][0] ), .B(
        \u_div/PartRem[60][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/SumTmp[58][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_59_1  ( .A(\u_div/PartRem[61][0] ), .B(
        \u_div/PartRem[61][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_1_3  ( .A(\u_div/PartRem[2][3] ), .B(
        \u_div/SumTmp[1][3] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_3  ( .A(\u_div/PartRem[3][3] ), .B(
        \u_div/SumTmp[2][3] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_3  ( .A(\u_div/PartRem[5][3] ), .B(
        \u_div/SumTmp[4][3] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_3  ( .A(\u_div/PartRem[7][3] ), .B(
        \u_div/SumTmp[6][3] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_9_3  ( .A(\u_div/PartRem[10][3] ), .B(
        \u_div/SumTmp[9][3] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_3  ( .A(\u_div/PartRem[12][3] ), .B(
        \u_div/SumTmp[11][3] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_3  ( .A(\u_div/PartRem[13][3] ), .B(
        \u_div/SumTmp[12][3] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_3  ( .A(\u_div/PartRem[15][3] ), .B(
        \u_div/SumTmp[14][3] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_3  ( .A(\u_div/PartRem[17][3] ), .B(
        \u_div/SumTmp[16][3] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_3  ( .A(\u_div/PartRem[18][3] ), .B(
        \u_div/SumTmp[17][3] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_3  ( .A(\u_div/PartRem[20][3] ), .B(
        \u_div/SumTmp[19][3] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_3  ( .A(\u_div/PartRem[22][3] ), .B(
        \u_div/SumTmp[21][3] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_3  ( .A(\u_div/PartRem[23][3] ), .B(
        \u_div/SumTmp[22][3] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_3  ( .A(\u_div/PartRem[25][3] ), .B(
        \u_div/SumTmp[24][3] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_3  ( .A(\u_div/PartRem[27][3] ), .B(
        \u_div/SumTmp[26][3] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_3  ( .A(\u_div/PartRem[28][3] ), .B(
        \u_div/SumTmp[27][3] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_3  ( .A(\u_div/PartRem[30][3] ), .B(
        \u_div/SumTmp[29][3] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_3  ( .A(\u_div/PartRem[32][3] ), .B(
        \u_div/SumTmp[31][3] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_3  ( .A(\u_div/PartRem[33][3] ), .B(
        \u_div/SumTmp[32][3] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_3  ( .A(\u_div/PartRem[35][3] ), .B(
        \u_div/SumTmp[34][3] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_3  ( .A(\u_div/PartRem[37][3] ), .B(
        \u_div/SumTmp[36][3] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_3  ( .A(\u_div/PartRem[38][3] ), .B(
        \u_div/SumTmp[37][3] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_3  ( .A(\u_div/PartRem[40][3] ), .B(
        \u_div/SumTmp[39][3] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_3  ( .A(\u_div/PartRem[42][3] ), .B(
        \u_div/SumTmp[41][3] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_3  ( .A(\u_div/PartRem[43][3] ), .B(
        \u_div/SumTmp[42][3] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_3  ( .A(\u_div/PartRem[45][3] ), .B(
        \u_div/SumTmp[44][3] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_3  ( .A(\u_div/PartRem[47][3] ), .B(
        \u_div/SumTmp[46][3] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_3  ( .A(\u_div/PartRem[48][3] ), .B(
        \u_div/SumTmp[47][3] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_3  ( .A(\u_div/PartRem[50][3] ), .B(
        \u_div/SumTmp[49][3] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_3  ( .A(\u_div/PartRem[52][3] ), .B(
        \u_div/SumTmp[51][3] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_3  ( .A(\u_div/PartRem[53][3] ), .B(
        \u_div/SumTmp[52][3] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_3  ( .A(\u_div/PartRem[55][3] ), .B(
        \u_div/SumTmp[54][3] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_3  ( .A(\u_div/PartRem[57][3] ), .B(
        \u_div/SumTmp[56][3] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_3  ( .A(\u_div/PartRem[58][3] ), .B(
        \u_div/SumTmp[57][3] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_3  ( .A(\u_div/PartRem[59][3] ), .B(
        \u_div/SumTmp[58][3] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_3  ( .A(\u_div/PartRem[63][0] ), .B(
        \u_div/SumTmp[59][3] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_3  ( .A(\u_div/PartRem[4][3] ), .B(
        \u_div/SumTmp[3][3] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_8_3  ( .A(\u_div/PartRem[9][3] ), .B(
        \u_div/SumTmp[8][3] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_3  ( .A(\u_div/PartRem[14][3] ), .B(
        \u_div/SumTmp[13][3] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_3  ( .A(\u_div/PartRem[19][3] ), .B(
        \u_div/SumTmp[18][3] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_3  ( .A(\u_div/PartRem[24][3] ), .B(
        \u_div/SumTmp[23][3] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_3  ( .A(\u_div/PartRem[29][3] ), .B(
        \u_div/SumTmp[28][3] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_3  ( .A(\u_div/PartRem[34][3] ), .B(
        \u_div/SumTmp[33][3] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_3  ( .A(\u_div/PartRem[39][3] ), .B(
        \u_div/SumTmp[38][3] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_3  ( .A(\u_div/PartRem[44][3] ), .B(
        \u_div/SumTmp[43][3] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_3  ( .A(\u_div/PartRem[49][3] ), .B(
        \u_div/SumTmp[48][3] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_3  ( .A(\u_div/PartRem[54][3] ), .B(
        \u_div/SumTmp[53][3] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/SumTmp[1][2] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][3] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_4  ( .A(\u_div/PartRem[64][0] ), .B(
        \u_div/SumTmp[59][4] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_3_1  ( .A(\u_div/SumTmp[3][1] ), .B(
        \u_div/SumTmp[3][1] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_4_1  ( .A(\u_div/SumTmp[4][1] ), .B(
        \u_div/SumTmp[4][1] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_0  ( .A(\u_div/PartRem[6][0] ), .B(
        \u_div/PartRem[6][0] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/SumTmp[4][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_13_1  ( .A(\u_div/SumTmp[13][1] ), .B(
        \u_div/SumTmp[13][1] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_18_1  ( .A(\u_div/SumTmp[18][1] ), .B(
        \u_div/SumTmp[18][1] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_23_1  ( .A(\u_div/SumTmp[23][1] ), .B(
        \u_div/SumTmp[23][1] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_0  ( .A(\u_div/PartRem[11][0] ), .B(
        \u_div/PartRem[11][0] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/SumTmp[9][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_14_1  ( .A(\u_div/SumTmp[14][1] ), .B(
        \u_div/SumTmp[14][1] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_0  ( .A(\u_div/PartRem[16][0] ), .B(
        \u_div/PartRem[16][0] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/SumTmp[14][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_0  ( .A(\u_div/PartRem[21][0] ), .B(
        \u_div/PartRem[21][0] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/SumTmp[19][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_24_1  ( .A(\u_div/SumTmp[24][1] ), .B(
        \u_div/SumTmp[24][1] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_0  ( .A(\u_div/PartRem[26][0] ), .B(
        \u_div/PartRem[26][0] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/SumTmp[24][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_12_1  ( .A(\u_div/SumTmp[12][1] ), .B(
        \u_div/SumTmp[12][1] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_17_1  ( .A(\u_div/SumTmp[17][1] ), .B(
        \u_div/SumTmp[17][1] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_22_1  ( .A(\u_div/SumTmp[22][1] ), .B(
        \u_div/SumTmp[22][1] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_6_1  ( .A(\u_div/SumTmp[6][1] ), .B(
        \u_div/SumTmp[6][1] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_11_1  ( .A(\u_div/SumTmp[11][1] ), .B(
        \u_div/SumTmp[11][1] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_16_1  ( .A(\u_div/SumTmp[16][1] ), .B(
        \u_div/SumTmp[16][1] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_21_1  ( .A(\u_div/SumTmp[21][1] ), .B(
        \u_div/SumTmp[21][1] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_26_1  ( .A(\u_div/SumTmp[26][1] ), .B(
        \u_div/SumTmp[26][1] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_27_1  ( .A(\u_div/SumTmp[27][1] ), .B(
        \u_div/SumTmp[27][1] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_29_1  ( .A(\u_div/SumTmp[29][1] ), .B(
        \u_div/SumTmp[29][1] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_0  ( .A(\u_div/PartRem[31][0] ), .B(
        \u_div/PartRem[31][0] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/SumTmp[29][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_31_1  ( .A(\u_div/SumTmp[31][1] ), .B(
        \u_div/SumTmp[31][1] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_32_1  ( .A(\u_div/SumTmp[32][1] ), .B(
        \u_div/SumTmp[32][1] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_33_1  ( .A(\u_div/SumTmp[33][1] ), .B(
        \u_div/SumTmp[33][1] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_34_1  ( .A(\u_div/SumTmp[34][1] ), .B(
        \u_div/SumTmp[34][1] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_0  ( .A(\u_div/PartRem[36][0] ), .B(
        \u_div/PartRem[36][0] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/SumTmp[34][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_36_1  ( .A(\u_div/SumTmp[36][1] ), .B(
        \u_div/SumTmp[36][1] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_37_1  ( .A(\u_div/SumTmp[37][1] ), .B(
        \u_div/SumTmp[37][1] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_39_1  ( .A(\u_div/SumTmp[39][1] ), .B(
        \u_div/SumTmp[39][1] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_0  ( .A(\u_div/PartRem[41][0] ), .B(
        \u_div/PartRem[41][0] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/SumTmp[39][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_41_1  ( .A(\u_div/SumTmp[41][1] ), .B(
        \u_div/SumTmp[41][1] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_42_1  ( .A(\u_div/SumTmp[42][1] ), .B(
        \u_div/SumTmp[42][1] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_43_1  ( .A(\u_div/SumTmp[43][1] ), .B(
        \u_div/SumTmp[43][1] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_44_1  ( .A(\u_div/SumTmp[44][1] ), .B(
        \u_div/SumTmp[44][1] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_0  ( .A(\u_div/PartRem[46][0] ), .B(
        \u_div/PartRem[46][0] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/SumTmp[44][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_46_1  ( .A(\u_div/SumTmp[46][1] ), .B(
        \u_div/SumTmp[46][1] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_47_1  ( .A(\u_div/SumTmp[47][1] ), .B(
        \u_div/SumTmp[47][1] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_0  ( .A(\u_div/PartRem[51][0] ), .B(
        \u_div/PartRem[51][0] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/SumTmp[49][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_51_1  ( .A(\u_div/SumTmp[51][1] ), .B(
        \u_div/SumTmp[51][1] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_52_1  ( .A(\u_div/SumTmp[52][1] ), .B(
        \u_div/SumTmp[52][1] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_53_1  ( .A(\u_div/SumTmp[53][1] ), .B(
        \u_div/SumTmp[53][1] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_54_1  ( .A(\u_div/SumTmp[54][1] ), .B(
        \u_div/SumTmp[54][1] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_0  ( .A(\u_div/PartRem[56][0] ), .B(
        \u_div/PartRem[56][0] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/SumTmp[54][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_57_1  ( .A(\u_div/SumTmp[57][1] ), .B(
        \u_div/SumTmp[57][1] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_58_1  ( .A(\u_div/SumTmp[58][1] ), .B(
        \u_div/SumTmp[58][1] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_2_1  ( .A(\u_div/SumTmp[2][1] ), .B(
        \u_div/SumTmp[2][1] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_3  ( .A(\u_div/PartRem[6][3] ), .B(
        \u_div/SumTmp[5][3] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_3  ( .A(\u_div/PartRem[11][3] ), .B(
        \u_div/SumTmp[10][3] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_3  ( .A(\u_div/PartRem[16][3] ), .B(
        \u_div/SumTmp[15][3] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_3  ( .A(\u_div/PartRem[21][3] ), .B(
        \u_div/SumTmp[20][3] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_3  ( .A(\u_div/PartRem[26][3] ), .B(
        \u_div/SumTmp[25][3] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_3  ( .A(\u_div/PartRem[31][3] ), .B(
        \u_div/SumTmp[30][3] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_3  ( .A(\u_div/PartRem[36][3] ), .B(
        \u_div/SumTmp[35][3] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_3  ( .A(\u_div/PartRem[41][3] ), .B(
        \u_div/SumTmp[40][3] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_3  ( .A(\u_div/PartRem[46][3] ), .B(
        \u_div/SumTmp[45][3] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_3  ( .A(\u_div/PartRem[51][3] ), .B(
        \u_div/SumTmp[50][3] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_3  ( .A(\u_div/PartRem[56][3] ), .B(
        \u_div/SumTmp[55][3] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_1_4  ( .A(\u_div/PartRem[2][4] ), .B(
        \u_div/SumTmp[1][4] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_4  ( .A(\u_div/PartRem[7][4] ), .B(
        \u_div/SumTmp[6][4] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_4  ( .A(\u_div/PartRem[12][4] ), .B(
        \u_div/SumTmp[11][4] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_4  ( .A(\u_div/PartRem[17][4] ), .B(
        \u_div/SumTmp[16][4] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_4  ( .A(\u_div/PartRem[22][4] ), .B(
        \u_div/SumTmp[21][4] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_4  ( .A(\u_div/PartRem[27][4] ), .B(
        \u_div/SumTmp[26][4] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_4  ( .A(\u_div/PartRem[32][4] ), .B(
        \u_div/SumTmp[31][4] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_4  ( .A(\u_div/PartRem[37][4] ), .B(
        \u_div/SumTmp[36][4] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_4  ( .A(\u_div/PartRem[42][4] ), .B(
        \u_div/SumTmp[41][4] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_4  ( .A(\u_div/PartRem[47][4] ), .B(
        \u_div/SumTmp[46][4] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_4  ( .A(\u_div/PartRem[52][4] ), .B(
        \u_div/SumTmp[51][4] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_4  ( .A(\u_div/PartRem[3][4] ), .B(
        \u_div/SumTmp[2][4] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_4  ( .A(\u_div/PartRem[4][4] ), .B(
        \u_div/SumTmp[3][4] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_4  ( .A(\u_div/PartRem[5][4] ), .B(
        \u_div/SumTmp[4][4] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_4  ( .A(\u_div/PartRem[6][4] ), .B(
        \u_div/SumTmp[5][4] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_4  ( .A(\u_div/PartRem[8][4] ), .B(
        \u_div/SumTmp[7][4] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_4  ( .A(\u_div/PartRem[15][4] ), .B(
        \u_div/SumTmp[14][4] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_4  ( .A(\u_div/PartRem[14][4] ), .B(
        \u_div/SumTmp[13][4] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_4  ( .A(\u_div/PartRem[19][4] ), .B(
        \u_div/SumTmp[18][4] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_4  ( .A(\u_div/PartRem[13][4] ), .B(
        \u_div/SumTmp[12][4] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_4  ( .A(\u_div/PartRem[18][4] ), .B(
        \u_div/SumTmp[17][4] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_4  ( .A(\u_div/PartRem[23][4] ), .B(
        \u_div/SumTmp[22][4] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_4  ( .A(\u_div/PartRem[24][4] ), .B(
        \u_div/SumTmp[23][4] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_4  ( .A(\u_div/PartRem[11][4] ), .B(
        \u_div/SumTmp[10][4] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_4  ( .A(\u_div/PartRem[16][4] ), .B(
        \u_div/SumTmp[15][4] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_4  ( .A(\u_div/PartRem[21][4] ), .B(
        \u_div/SumTmp[20][4] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_4  ( .A(\u_div/PartRem[26][4] ), .B(
        \u_div/SumTmp[25][4] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_4  ( .A(\u_div/PartRem[25][4] ), .B(
        \u_div/SumTmp[24][4] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_4  ( .A(\u_div/PartRem[28][4] ), .B(
        \u_div/SumTmp[27][4] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_4  ( .A(\u_div/PartRem[30][4] ), .B(
        \u_div/SumTmp[29][4] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_4  ( .A(\u_div/PartRem[31][4] ), .B(
        \u_div/SumTmp[30][4] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_4  ( .A(\u_div/PartRem[34][4] ), .B(
        \u_div/SumTmp[33][4] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_4  ( .A(\u_div/PartRem[33][4] ), .B(
        \u_div/SumTmp[32][4] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_4  ( .A(\u_div/PartRem[35][4] ), .B(
        \u_div/SumTmp[34][4] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_4  ( .A(\u_div/PartRem[36][4] ), .B(
        \u_div/SumTmp[35][4] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_4  ( .A(\u_div/PartRem[38][4] ), .B(
        \u_div/SumTmp[37][4] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_4  ( .A(\u_div/PartRem[40][4] ), .B(
        \u_div/SumTmp[39][4] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_4  ( .A(\u_div/PartRem[41][4] ), .B(
        \u_div/SumTmp[40][4] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_4  ( .A(\u_div/PartRem[44][4] ), .B(
        \u_div/SumTmp[43][4] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_4  ( .A(\u_div/PartRem[43][4] ), .B(
        \u_div/SumTmp[42][4] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_4  ( .A(\u_div/PartRem[45][4] ), .B(
        \u_div/SumTmp[44][4] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_4  ( .A(\u_div/PartRem[46][4] ), .B(
        \u_div/SumTmp[45][4] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_4  ( .A(\u_div/PartRem[48][4] ), .B(
        \u_div/SumTmp[47][4] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_4  ( .A(\u_div/PartRem[51][4] ), .B(
        \u_div/SumTmp[50][4] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_4  ( .A(\u_div/PartRem[55][4] ), .B(
        \u_div/SumTmp[54][4] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_4  ( .A(\u_div/PartRem[53][4] ), .B(
        \u_div/SumTmp[52][4] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_4  ( .A(\u_div/PartRem[54][4] ), .B(
        \u_div/SumTmp[53][4] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_4  ( .A(\u_div/PartRem[58][4] ), .B(
        \u_div/SumTmp[57][4] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_4  ( .A(\u_div/PartRem[56][4] ), .B(
        \u_div/SumTmp[55][4] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_4  ( .A(\u_div/PartRem[59][4] ), .B(
        \u_div/SumTmp[58][4] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_8_4  ( .A(\u_div/PartRem[9][4] ), .B(
        \u_div/SumTmp[8][4] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][5] ) );
  CLKMX2X6 \u_div/u_mx_PartRem_1_8_1  ( .A(\u_div/SumTmp[8][1] ), .B(
        \u_div/SumTmp[8][1] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_8_0  ( .A(\u_div/PartRem[9][0] ), .B(
        \u_div/PartRem[9][0] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/SumTmp[7][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_9_4  ( .A(\u_div/PartRem[10][4] ), .B(
        \u_div/SumTmp[9][4] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][5] ) );
  MX2X6 \u_div/u_mx_PartRem_1_9_1  ( .A(\u_div/SumTmp[9][1] ), .B(
        \u_div/SumTmp[9][1] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_9_0  ( .A(\u_div/PartRem[10][0] ), .B(
        \u_div/PartRem[10][0] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/SumTmp[8][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_19_4  ( .A(\u_div/PartRem[20][4] ), .B(
        \u_div/SumTmp[19][4] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][5] ) );
  MX2X6 \u_div/u_mx_PartRem_1_19_1  ( .A(\u_div/SumTmp[19][1] ), .B(
        \u_div/SumTmp[19][1] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_19_0  ( .A(\u_div/PartRem[20][0] ), .B(
        \u_div/PartRem[20][0] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/SumTmp[18][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_28_4  ( .A(\u_div/PartRem[29][4] ), .B(
        \u_div/SumTmp[28][4] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][5] ) );
  CLKMX2X6 \u_div/u_mx_PartRem_1_28_1  ( .A(\u_div/SumTmp[28][1] ), .B(
        \u_div/SumTmp[28][1] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_28_0  ( .A(\u_div/PartRem[29][0] ), .B(
        \u_div/PartRem[29][0] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/SumTmp[27][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_38_4  ( .A(\u_div/PartRem[39][4] ), .B(
        \u_div/SumTmp[38][4] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][5] ) );
  CLKMX2X6 \u_div/u_mx_PartRem_1_38_1  ( .A(\u_div/SumTmp[38][1] ), .B(
        \u_div/SumTmp[38][1] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_38_0  ( .A(\u_div/PartRem[39][0] ), .B(
        \u_div/PartRem[39][0] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/SumTmp[37][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_48_4  ( .A(\u_div/PartRem[49][4] ), .B(
        \u_div/SumTmp[48][4] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][5] ) );
  CLKMX2X6 \u_div/u_mx_PartRem_1_48_1  ( .A(\u_div/SumTmp[48][1] ), .B(
        \u_div/SumTmp[48][1] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_48_0  ( .A(\u_div/PartRem[49][0] ), .B(
        \u_div/PartRem[49][0] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/SumTmp[47][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_49_4  ( .A(\u_div/PartRem[50][4] ), .B(
        \u_div/SumTmp[49][4] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][5] ) );
  MX2X6 \u_div/u_mx_PartRem_1_49_1  ( .A(\u_div/SumTmp[49][1] ), .B(
        \u_div/SumTmp[49][1] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_49_0  ( .A(\u_div/PartRem[50][0] ), .B(
        \u_div/PartRem[50][0] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/SumTmp[48][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_56_4  ( .A(\u_div/PartRem[57][4] ), .B(
        \u_div/SumTmp[56][4] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][5] ) );
  CLKMX2X6 \u_div/u_mx_PartRem_1_56_1  ( .A(\u_div/SumTmp[56][1] ), .B(
        \u_div/SumTmp[56][1] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][2] ) );
  CLKMX2X4 \u_div/u_mx_PartRem_1_56_0  ( .A(\u_div/PartRem[57][0] ), .B(
        \u_div/PartRem[57][0] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/SumTmp[55][1] ) );
  MX2X6 \u_div/u_mx_PartRem_1_7_1  ( .A(\u_div/SumTmp[7][1] ), .B(
        \u_div/SumTmp[7][1] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][2] ) );
  MX2X4 \u_div/u_mx_PartRem_1_7_3  ( .A(\u_div/PartRem[8][3] ), .B(
        \u_div/SumTmp[7][3] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][4] ) );
  OR2X2 U1 ( .A(\u_div/PartRem[11][5] ), .B(\u_div/u_add_PartRem_2_10/n2 ), 
        .Y(\u_div/CryTmp[10][6] ) );
  MXI2X4 U2 ( .A(\u_div/SumTmp[7][2] ), .B(\u_div/PartRem[8][2] ), .S0(
        \u_div/CryTmp[7][6] ), .Y(\u_div/PartRem[7][3] ) );
  OR2X6 U3 ( .A(\u_div/PartRem[8][5] ), .B(\u_div/u_add_PartRem_2_7/n2 ), .Y(
        \u_div/CryTmp[7][6] ) );
  OR2X8 U4 ( .A(\u_div/PartRem[7][5] ), .B(\u_div/u_add_PartRem_2_6/n2 ), .Y(
        \u_div/CryTmp[6][6] ) );
  ADDHX2 U5 ( .A(\u_div/PartRem[7][4] ), .B(\u_div/u_add_PartRem_2_6/n3 ), 
        .CO(\u_div/u_add_PartRem_2_6/n2 ), .S(\u_div/SumTmp[6][4] ) );
  OR2X8 U6 ( .A(\u_div/PartRem[6][5] ), .B(\u_div/u_add_PartRem_2_5/n2 ), .Y(
        \u_div/CryTmp[5][6] ) );
  ADDHX2 U7 ( .A(\u_div/PartRem[6][4] ), .B(\u_div/u_add_PartRem_2_5/n3 ), 
        .CO(\u_div/u_add_PartRem_2_5/n2 ), .S(\u_div/SumTmp[5][4] ) );
  OR2X8 U8 ( .A(\u_div/PartRem[5][5] ), .B(\u_div/u_add_PartRem_2_4/n2 ), .Y(
        \u_div/CryTmp[4][6] ) );
  ADDHX2 U9 ( .A(\u_div/PartRem[5][4] ), .B(\u_div/u_add_PartRem_2_4/n3 ), 
        .CO(\u_div/u_add_PartRem_2_4/n2 ), .S(\u_div/SumTmp[4][4] ) );
  OR2X8 U10 ( .A(\u_div/PartRem[4][5] ), .B(\u_div/u_add_PartRem_2_3/n2 ), .Y(
        \u_div/CryTmp[3][6] ) );
  ADDHX2 U11 ( .A(\u_div/PartRem[4][4] ), .B(\u_div/u_add_PartRem_2_3/n3 ), 
        .CO(\u_div/u_add_PartRem_2_3/n2 ), .S(\u_div/SumTmp[3][4] ) );
  OR2X8 U12 ( .A(\u_div/PartRem[3][5] ), .B(\u_div/u_add_PartRem_2_2/n2 ), .Y(
        \u_div/CryTmp[2][6] ) );
  ADDHX2 U13 ( .A(\u_div/PartRem[3][4] ), .B(\u_div/u_add_PartRem_2_2/n3 ), 
        .CO(\u_div/u_add_PartRem_2_2/n2 ), .S(\u_div/SumTmp[2][4] ) );
  OR2X8 U14 ( .A(\u_div/PartRem[59][5] ), .B(\u_div/u_add_PartRem_2_58/n2 ), 
        .Y(\u_div/CryTmp[58][6] ) );
  ADDHX2 U15 ( .A(\u_div/PartRem[59][4] ), .B(\u_div/u_add_PartRem_2_58/n3 ), 
        .CO(\u_div/u_add_PartRem_2_58/n2 ), .S(\u_div/SumTmp[58][4] ) );
  XOR2XL U16 ( .A(\u_div/CryTmp[56][6] ), .B(n3), .Y(\u_div/QInv[56] ) );
  MXI2X4 U17 ( .A(\u_div/SumTmp[56][2] ), .B(\u_div/PartRem[57][2] ), .S0(
        \u_div/CryTmp[56][6] ), .Y(\u_div/PartRem[56][3] ) );
  OR2X6 U18 ( .A(\u_div/PartRem[57][5] ), .B(\u_div/u_add_PartRem_2_56/n2 ), 
        .Y(\u_div/CryTmp[56][6] ) );
  XOR2XL U19 ( .A(\u_div/CryTmp[49][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[49] ) );
  MXI2X4 U20 ( .A(\u_div/SumTmp[49][2] ), .B(\u_div/PartRem[50][2] ), .S0(
        \u_div/CryTmp[49][6] ), .Y(\u_div/PartRem[49][3] ) );
  OR2X6 U21 ( .A(\u_div/PartRem[50][5] ), .B(\u_div/u_add_PartRem_2_49/n2 ), 
        .Y(\u_div/CryTmp[49][6] ) );
  XOR2XL U22 ( .A(\u_div/CryTmp[48][6] ), .B(n3), .Y(\u_div/QInv[48] ) );
  MXI2X4 U23 ( .A(\u_div/SumTmp[48][2] ), .B(\u_div/PartRem[49][2] ), .S0(
        \u_div/CryTmp[48][6] ), .Y(\u_div/PartRem[48][3] ) );
  OR2X6 U24 ( .A(\u_div/PartRem[49][5] ), .B(\u_div/u_add_PartRem_2_48/n2 ), 
        .Y(\u_div/CryTmp[48][6] ) );
  OR2X8 U25 ( .A(\u_div/PartRem[40][5] ), .B(\u_div/u_add_PartRem_2_39/n2 ), 
        .Y(\u_div/CryTmp[39][6] ) );
  ADDHX2 U26 ( .A(\u_div/PartRem[40][4] ), .B(\u_div/u_add_PartRem_2_39/n3 ), 
        .CO(\u_div/u_add_PartRem_2_39/n2 ), .S(\u_div/SumTmp[39][4] ) );
  XOR2XL U27 ( .A(\u_div/CryTmp[38][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[38] ) );
  MXI2X4 U28 ( .A(\u_div/SumTmp[38][2] ), .B(\u_div/PartRem[39][2] ), .S0(
        \u_div/CryTmp[38][6] ), .Y(\u_div/PartRem[38][3] ) );
  OR2X6 U29 ( .A(\u_div/PartRem[39][5] ), .B(\u_div/u_add_PartRem_2_38/n2 ), 
        .Y(\u_div/CryTmp[38][6] ) );
  OR2X8 U30 ( .A(\u_div/PartRem[30][5] ), .B(\u_div/u_add_PartRem_2_29/n2 ), 
        .Y(\u_div/CryTmp[29][6] ) );
  ADDHX2 U31 ( .A(\u_div/PartRem[30][4] ), .B(\u_div/u_add_PartRem_2_29/n3 ), 
        .CO(\u_div/u_add_PartRem_2_29/n2 ), .S(\u_div/SumTmp[29][4] ) );
  XOR2XL U32 ( .A(\u_div/CryTmp[28][6] ), .B(n5), .Y(\u_div/QInv[28] ) );
  MXI2X4 U33 ( .A(\u_div/SumTmp[28][2] ), .B(\u_div/PartRem[29][2] ), .S0(
        \u_div/CryTmp[28][6] ), .Y(\u_div/PartRem[28][3] ) );
  OR2X6 U34 ( .A(\u_div/PartRem[29][5] ), .B(\u_div/u_add_PartRem_2_28/n2 ), 
        .Y(\u_div/CryTmp[28][6] ) );
  XOR2XL U35 ( .A(\u_div/CryTmp[19][6] ), .B(n3), .Y(\u_div/QInv[19] ) );
  MXI2X4 U36 ( .A(\u_div/SumTmp[19][2] ), .B(\u_div/PartRem[20][2] ), .S0(
        \u_div/CryTmp[19][6] ), .Y(\u_div/PartRem[19][3] ) );
  OR2X6 U37 ( .A(\u_div/PartRem[20][5] ), .B(\u_div/u_add_PartRem_2_19/n2 ), 
        .Y(\u_div/CryTmp[19][6] ) );
  OR2X8 U38 ( .A(\u_div/PartRem[19][5] ), .B(\u_div/u_add_PartRem_2_18/n2 ), 
        .Y(\u_div/CryTmp[18][6] ) );
  ADDHX2 U39 ( .A(\u_div/PartRem[19][4] ), .B(\u_div/u_add_PartRem_2_18/n3 ), 
        .CO(\u_div/u_add_PartRem_2_18/n2 ), .S(\u_div/SumTmp[18][4] ) );
  XOR2XL U40 ( .A(\u_div/CryTmp[9][6] ), .B(n3), .Y(\u_div/QInv[9] ) );
  MXI2X4 U41 ( .A(\u_div/SumTmp[9][2] ), .B(\u_div/PartRem[10][2] ), .S0(
        \u_div/CryTmp[9][6] ), .Y(\u_div/PartRem[9][3] ) );
  OR2X6 U42 ( .A(\u_div/PartRem[10][5] ), .B(\u_div/u_add_PartRem_2_9/n2 ), 
        .Y(\u_div/CryTmp[9][6] ) );
  XOR2XL U43 ( .A(\u_div/CryTmp[8][6] ), .B(n3), .Y(\u_div/QInv[8] ) );
  MXI2X4 U44 ( .A(\u_div/SumTmp[8][2] ), .B(\u_div/PartRem[9][2] ), .S0(
        \u_div/CryTmp[8][6] ), .Y(\u_div/PartRem[8][3] ) );
  OR2X6 U45 ( .A(\u_div/PartRem[9][5] ), .B(\u_div/u_add_PartRem_2_8/n2 ), .Y(
        \u_div/CryTmp[8][6] ) );
  MXI2X1 U46 ( .A(\u_div/SumTmp[13][2] ), .B(\u_div/PartRem[14][2] ), .S0(
        \u_div/CryTmp[13][6] ), .Y(\u_div/PartRem[13][3] ) );
  MXI2X1 U47 ( .A(\u_div/SumTmp[18][2] ), .B(\u_div/PartRem[19][2] ), .S0(
        \u_div/CryTmp[18][6] ), .Y(\u_div/PartRem[18][3] ) );
  MXI2X1 U48 ( .A(\u_div/SumTmp[23][2] ), .B(\u_div/PartRem[24][2] ), .S0(
        \u_div/CryTmp[23][6] ), .Y(\u_div/PartRem[23][3] ) );
  MXI2X1 U49 ( .A(\u_div/SumTmp[33][2] ), .B(\u_div/PartRem[34][2] ), .S0(
        \u_div/CryTmp[33][6] ), .Y(\u_div/PartRem[33][3] ) );
  MXI2X1 U50 ( .A(\u_div/SumTmp[43][2] ), .B(\u_div/PartRem[44][2] ), .S0(
        \u_div/CryTmp[43][6] ), .Y(\u_div/PartRem[43][3] ) );
  MXI2X1 U51 ( .A(\u_div/SumTmp[53][2] ), .B(\u_div/PartRem[54][2] ), .S0(
        \u_div/CryTmp[53][6] ), .Y(\u_div/PartRem[53][3] ) );
  ADDHXL U52 ( .A(\u_div/PartRem[13][4] ), .B(\u_div/u_add_PartRem_2_12/n3 ), 
        .CO(\u_div/u_add_PartRem_2_12/n2 ), .S(\u_div/SumTmp[12][4] ) );
  ADDHXL U53 ( .A(\u_div/PartRem[12][4] ), .B(\u_div/u_add_PartRem_2_11/n3 ), 
        .CO(\u_div/u_add_PartRem_2_11/n2 ), .S(\u_div/SumTmp[11][4] ) );
  OR2X1 U54 ( .A(\u_div/PartRem[12][2] ), .B(\u_div/PartRem[12][3] ), .Y(
        \u_div/u_add_PartRem_2_11/n3 ) );
  ADDHXL U55 ( .A(\u_div/PartRem[15][4] ), .B(\u_div/u_add_PartRem_2_14/n3 ), 
        .CO(\u_div/u_add_PartRem_2_14/n2 ), .S(\u_div/SumTmp[14][4] ) );
  OR2X1 U56 ( .A(\u_div/PartRem[15][2] ), .B(\u_div/PartRem[15][3] ), .Y(
        \u_div/u_add_PartRem_2_14/n3 ) );
  ADDHXL U57 ( .A(\u_div/PartRem[14][4] ), .B(\u_div/u_add_PartRem_2_13/n3 ), 
        .CO(\u_div/u_add_PartRem_2_13/n2 ), .S(\u_div/SumTmp[13][4] ) );
  OR2X1 U58 ( .A(\u_div/PartRem[14][2] ), .B(\u_div/PartRem[14][3] ), .Y(
        \u_div/u_add_PartRem_2_13/n3 ) );
  ADDHXL U59 ( .A(\u_div/PartRem[16][4] ), .B(\u_div/u_add_PartRem_2_15/n3 ), 
        .CO(\u_div/u_add_PartRem_2_15/n2 ), .S(\u_div/SumTmp[15][4] ) );
  OR2X1 U60 ( .A(\u_div/PartRem[16][2] ), .B(\u_div/PartRem[16][3] ), .Y(
        \u_div/u_add_PartRem_2_15/n3 ) );
  ADDHXL U61 ( .A(\u_div/PartRem[17][4] ), .B(\u_div/u_add_PartRem_2_16/n3 ), 
        .CO(\u_div/u_add_PartRem_2_16/n2 ), .S(\u_div/SumTmp[16][4] ) );
  OR2X1 U62 ( .A(\u_div/PartRem[17][2] ), .B(\u_div/PartRem[17][3] ), .Y(
        \u_div/u_add_PartRem_2_16/n3 ) );
  ADDHXL U63 ( .A(\u_div/PartRem[18][4] ), .B(\u_div/u_add_PartRem_2_17/n3 ), 
        .CO(\u_div/u_add_PartRem_2_17/n2 ), .S(\u_div/SumTmp[17][4] ) );
  OR2X1 U64 ( .A(\u_div/PartRem[19][2] ), .B(\u_div/PartRem[19][3] ), .Y(
        \u_div/u_add_PartRem_2_18/n3 ) );
  ADDHXL U65 ( .A(\u_div/PartRem[20][4] ), .B(\u_div/u_add_PartRem_2_19/n3 ), 
        .CO(\u_div/u_add_PartRem_2_19/n2 ), .S(\u_div/SumTmp[19][4] ) );
  OR2X1 U66 ( .A(\u_div/PartRem[20][2] ), .B(\u_div/PartRem[20][3] ), .Y(
        \u_div/u_add_PartRem_2_19/n3 ) );
  ADDHXL U67 ( .A(\u_div/PartRem[24][4] ), .B(\u_div/u_add_PartRem_2_23/n3 ), 
        .CO(\u_div/u_add_PartRem_2_23/n2 ), .S(\u_div/SumTmp[23][4] ) );
  OR2X1 U68 ( .A(\u_div/PartRem[24][2] ), .B(\u_div/PartRem[24][3] ), .Y(
        \u_div/u_add_PartRem_2_23/n3 ) );
  ADDHXL U69 ( .A(\u_div/PartRem[23][4] ), .B(\u_div/u_add_PartRem_2_22/n3 ), 
        .CO(\u_div/u_add_PartRem_2_22/n2 ), .S(\u_div/SumTmp[22][4] ) );
  ADDHXL U70 ( .A(\u_div/PartRem[22][4] ), .B(\u_div/u_add_PartRem_2_21/n3 ), 
        .CO(\u_div/u_add_PartRem_2_21/n2 ), .S(\u_div/SumTmp[21][4] ) );
  OR2X1 U71 ( .A(\u_div/PartRem[22][2] ), .B(\u_div/PartRem[22][3] ), .Y(
        \u_div/u_add_PartRem_2_21/n3 ) );
  ADDHXL U72 ( .A(\u_div/PartRem[21][4] ), .B(\u_div/u_add_PartRem_2_20/n3 ), 
        .CO(\u_div/u_add_PartRem_2_20/n2 ), .S(\u_div/SumTmp[20][4] ) );
  OR2X1 U73 ( .A(\u_div/PartRem[21][2] ), .B(\u_div/PartRem[21][3] ), .Y(
        \u_div/u_add_PartRem_2_20/n3 ) );
  MXI2X1 U74 ( .A(\u_div/SumTmp[3][2] ), .B(\u_div/PartRem[4][2] ), .S0(
        \u_div/CryTmp[3][6] ), .Y(\u_div/PartRem[3][3] ) );
  OR2X1 U75 ( .A(\u_div/PartRem[7][2] ), .B(\u_div/PartRem[7][3] ), .Y(
        \u_div/u_add_PartRem_2_6/n3 ) );
  ADDHXL U76 ( .A(\u_div/PartRem[11][4] ), .B(\u_div/u_add_PartRem_2_10/n3 ), 
        .CO(\u_div/u_add_PartRem_2_10/n2 ), .S(\u_div/SumTmp[10][4] ) );
  OR2X1 U77 ( .A(\u_div/PartRem[11][2] ), .B(\u_div/PartRem[11][3] ), .Y(
        \u_div/u_add_PartRem_2_10/n3 ) );
  OR2X1 U78 ( .A(\u_div/PartRem[4][2] ), .B(\u_div/PartRem[4][3] ), .Y(
        \u_div/u_add_PartRem_2_3/n3 ) );
  ADDHXL U79 ( .A(\u_div/PartRem[8][4] ), .B(\u_div/u_add_PartRem_2_7/n3 ), 
        .CO(\u_div/u_add_PartRem_2_7/n2 ), .S(\u_div/SumTmp[7][4] ) );
  ADDHXL U80 ( .A(\u_div/PartRem[10][4] ), .B(\u_div/u_add_PartRem_2_9/n3 ), 
        .CO(\u_div/u_add_PartRem_2_9/n2 ), .S(\u_div/SumTmp[9][4] ) );
  OR2X1 U81 ( .A(\u_div/PartRem[10][2] ), .B(\u_div/PartRem[10][3] ), .Y(
        \u_div/u_add_PartRem_2_9/n3 ) );
  ADDHXL U82 ( .A(\u_div/PartRem[9][4] ), .B(\u_div/u_add_PartRem_2_8/n3 ), 
        .CO(\u_div/u_add_PartRem_2_8/n2 ), .S(\u_div/SumTmp[8][4] ) );
  OR2X1 U83 ( .A(\u_div/PartRem[9][2] ), .B(\u_div/PartRem[9][3] ), .Y(
        \u_div/u_add_PartRem_2_8/n3 ) );
  OR2X1 U84 ( .A(\u_div/PartRem[6][2] ), .B(\u_div/PartRem[6][3] ), .Y(
        \u_div/u_add_PartRem_2_5/n3 ) );
  OR2X1 U85 ( .A(\u_div/PartRem[5][2] ), .B(\u_div/PartRem[5][3] ), .Y(
        \u_div/u_add_PartRem_2_4/n3 ) );
  ADDHXL U86 ( .A(\u_div/PartRem[25][4] ), .B(\u_div/u_add_PartRem_2_24/n3 ), 
        .CO(\u_div/u_add_PartRem_2_24/n2 ), .S(\u_div/SumTmp[24][4] ) );
  OR2X1 U87 ( .A(\u_div/PartRem[25][2] ), .B(\u_div/PartRem[25][3] ), .Y(
        \u_div/u_add_PartRem_2_24/n3 ) );
  ADDHXL U88 ( .A(\u_div/PartRem[26][4] ), .B(\u_div/u_add_PartRem_2_25/n3 ), 
        .CO(\u_div/u_add_PartRem_2_25/n2 ), .S(\u_div/SumTmp[25][4] ) );
  OR2X1 U89 ( .A(\u_div/PartRem[26][2] ), .B(\u_div/PartRem[26][3] ), .Y(
        \u_div/u_add_PartRem_2_25/n3 ) );
  ADDHXL U90 ( .A(\u_div/PartRem[27][4] ), .B(\u_div/u_add_PartRem_2_26/n3 ), 
        .CO(\u_div/u_add_PartRem_2_26/n2 ), .S(\u_div/SumTmp[26][4] ) );
  OR2X1 U91 ( .A(\u_div/PartRem[27][2] ), .B(\u_div/PartRem[27][3] ), .Y(
        \u_div/u_add_PartRem_2_26/n3 ) );
  ADDHXL U92 ( .A(\u_div/PartRem[28][4] ), .B(\u_div/u_add_PartRem_2_27/n3 ), 
        .CO(\u_div/u_add_PartRem_2_27/n2 ), .S(\u_div/SumTmp[27][4] ) );
  ADDHXL U93 ( .A(\u_div/PartRem[29][4] ), .B(\u_div/u_add_PartRem_2_28/n3 ), 
        .CO(\u_div/u_add_PartRem_2_28/n2 ), .S(\u_div/SumTmp[28][4] ) );
  OR2X1 U94 ( .A(\u_div/PartRem[29][2] ), .B(\u_div/PartRem[29][3] ), .Y(
        \u_div/u_add_PartRem_2_28/n3 ) );
  OR2X1 U95 ( .A(\u_div/PartRem[30][2] ), .B(\u_div/PartRem[30][3] ), .Y(
        \u_div/u_add_PartRem_2_29/n3 ) );
  ADDHXL U96 ( .A(\u_div/PartRem[31][4] ), .B(\u_div/u_add_PartRem_2_30/n3 ), 
        .CO(\u_div/u_add_PartRem_2_30/n2 ), .S(\u_div/SumTmp[30][4] ) );
  OR2X1 U97 ( .A(\u_div/PartRem[31][2] ), .B(\u_div/PartRem[31][3] ), .Y(
        \u_div/u_add_PartRem_2_30/n3 ) );
  ADDHXL U98 ( .A(\u_div/PartRem[33][4] ), .B(\u_div/u_add_PartRem_2_32/n3 ), 
        .CO(\u_div/u_add_PartRem_2_32/n2 ), .S(\u_div/SumTmp[32][4] ) );
  ADDHXL U99 ( .A(\u_div/PartRem[32][4] ), .B(\u_div/u_add_PartRem_2_31/n3 ), 
        .CO(\u_div/u_add_PartRem_2_31/n2 ), .S(\u_div/SumTmp[31][4] ) );
  OR2X1 U100 ( .A(\u_div/PartRem[32][2] ), .B(\u_div/PartRem[32][3] ), .Y(
        \u_div/u_add_PartRem_2_31/n3 ) );
  ADDHXL U101 ( .A(\u_div/PartRem[34][4] ), .B(\u_div/u_add_PartRem_2_33/n3 ), 
        .CO(\u_div/u_add_PartRem_2_33/n2 ), .S(\u_div/SumTmp[33][4] ) );
  OR2X1 U102 ( .A(\u_div/PartRem[34][2] ), .B(\u_div/PartRem[34][3] ), .Y(
        \u_div/u_add_PartRem_2_33/n3 ) );
  ADDHXL U103 ( .A(\u_div/PartRem[35][4] ), .B(\u_div/u_add_PartRem_2_34/n3 ), 
        .CO(\u_div/u_add_PartRem_2_34/n2 ), .S(\u_div/SumTmp[34][4] ) );
  OR2X1 U104 ( .A(\u_div/PartRem[35][2] ), .B(\u_div/PartRem[35][3] ), .Y(
        \u_div/u_add_PartRem_2_34/n3 ) );
  ADDHXL U105 ( .A(\u_div/PartRem[36][4] ), .B(\u_div/u_add_PartRem_2_35/n3 ), 
        .CO(\u_div/u_add_PartRem_2_35/n2 ), .S(\u_div/SumTmp[35][4] ) );
  OR2X1 U106 ( .A(\u_div/PartRem[36][2] ), .B(\u_div/PartRem[36][3] ), .Y(
        \u_div/u_add_PartRem_2_35/n3 ) );
  ADDHXL U107 ( .A(\u_div/PartRem[37][4] ), .B(\u_div/u_add_PartRem_2_36/n3 ), 
        .CO(\u_div/u_add_PartRem_2_36/n2 ), .S(\u_div/SumTmp[36][4] ) );
  OR2X1 U108 ( .A(\u_div/PartRem[37][2] ), .B(\u_div/PartRem[37][3] ), .Y(
        \u_div/u_add_PartRem_2_36/n3 ) );
  ADDHXL U109 ( .A(\u_div/PartRem[38][4] ), .B(\u_div/u_add_PartRem_2_37/n3 ), 
        .CO(\u_div/u_add_PartRem_2_37/n2 ), .S(\u_div/SumTmp[37][4] ) );
  ADDHXL U110 ( .A(\u_div/PartRem[39][4] ), .B(\u_div/u_add_PartRem_2_38/n3 ), 
        .CO(\u_div/u_add_PartRem_2_38/n2 ), .S(\u_div/SumTmp[38][4] ) );
  OR2X1 U111 ( .A(\u_div/PartRem[39][2] ), .B(\u_div/PartRem[39][3] ), .Y(
        \u_div/u_add_PartRem_2_38/n3 ) );
  OR2X1 U112 ( .A(\u_div/PartRem[40][2] ), .B(\u_div/PartRem[40][3] ), .Y(
        \u_div/u_add_PartRem_2_39/n3 ) );
  ADDHXL U113 ( .A(\u_div/PartRem[41][4] ), .B(\u_div/u_add_PartRem_2_40/n3 ), 
        .CO(\u_div/u_add_PartRem_2_40/n2 ), .S(\u_div/SumTmp[40][4] ) );
  OR2X1 U114 ( .A(\u_div/PartRem[41][2] ), .B(\u_div/PartRem[41][3] ), .Y(
        \u_div/u_add_PartRem_2_40/n3 ) );
  ADDHXL U115 ( .A(\u_div/PartRem[42][4] ), .B(\u_div/u_add_PartRem_2_41/n3 ), 
        .CO(\u_div/u_add_PartRem_2_41/n2 ), .S(\u_div/SumTmp[41][4] ) );
  OR2X1 U116 ( .A(\u_div/PartRem[42][2] ), .B(\u_div/PartRem[42][3] ), .Y(
        \u_div/u_add_PartRem_2_41/n3 ) );
  ADDHXL U117 ( .A(\u_div/PartRem[43][4] ), .B(\u_div/u_add_PartRem_2_42/n3 ), 
        .CO(\u_div/u_add_PartRem_2_42/n2 ), .S(\u_div/SumTmp[42][4] ) );
  ADDHXL U118 ( .A(\u_div/PartRem[44][4] ), .B(\u_div/u_add_PartRem_2_43/n3 ), 
        .CO(\u_div/u_add_PartRem_2_43/n2 ), .S(\u_div/SumTmp[43][4] ) );
  OR2X1 U119 ( .A(\u_div/PartRem[44][2] ), .B(\u_div/PartRem[44][3] ), .Y(
        \u_div/u_add_PartRem_2_43/n3 ) );
  ADDHXL U120 ( .A(\u_div/PartRem[45][4] ), .B(\u_div/u_add_PartRem_2_44/n3 ), 
        .CO(\u_div/u_add_PartRem_2_44/n2 ), .S(\u_div/SumTmp[44][4] ) );
  OR2X1 U121 ( .A(\u_div/PartRem[45][2] ), .B(\u_div/PartRem[45][3] ), .Y(
        \u_div/u_add_PartRem_2_44/n3 ) );
  ADDHXL U122 ( .A(\u_div/PartRem[46][4] ), .B(\u_div/u_add_PartRem_2_45/n3 ), 
        .CO(\u_div/u_add_PartRem_2_45/n2 ), .S(\u_div/SumTmp[45][4] ) );
  OR2X1 U123 ( .A(\u_div/PartRem[46][2] ), .B(\u_div/PartRem[46][3] ), .Y(
        \u_div/u_add_PartRem_2_45/n3 ) );
  ADDHXL U124 ( .A(\u_div/PartRem[47][4] ), .B(\u_div/u_add_PartRem_2_46/n3 ), 
        .CO(\u_div/u_add_PartRem_2_46/n2 ), .S(\u_div/SumTmp[46][4] ) );
  OR2X1 U125 ( .A(\u_div/PartRem[47][2] ), .B(\u_div/PartRem[47][3] ), .Y(
        \u_div/u_add_PartRem_2_46/n3 ) );
  ADDHXL U126 ( .A(\u_div/PartRem[48][4] ), .B(\u_div/u_add_PartRem_2_47/n3 ), 
        .CO(\u_div/u_add_PartRem_2_47/n2 ), .S(\u_div/SumTmp[47][4] ) );
  ADDHXL U127 ( .A(\u_div/PartRem[50][4] ), .B(\u_div/u_add_PartRem_2_49/n3 ), 
        .CO(\u_div/u_add_PartRem_2_49/n2 ), .S(\u_div/SumTmp[49][4] ) );
  OR2X1 U128 ( .A(\u_div/PartRem[50][2] ), .B(\u_div/PartRem[50][3] ), .Y(
        \u_div/u_add_PartRem_2_49/n3 ) );
  ADDHXL U129 ( .A(\u_div/PartRem[49][4] ), .B(\u_div/u_add_PartRem_2_48/n3 ), 
        .CO(\u_div/u_add_PartRem_2_48/n2 ), .S(\u_div/SumTmp[48][4] ) );
  OR2X1 U130 ( .A(\u_div/PartRem[49][2] ), .B(\u_div/PartRem[49][3] ), .Y(
        \u_div/u_add_PartRem_2_48/n3 ) );
  ADDHXL U131 ( .A(\u_div/PartRem[51][4] ), .B(\u_div/u_add_PartRem_2_50/n3 ), 
        .CO(\u_div/u_add_PartRem_2_50/n2 ), .S(\u_div/SumTmp[50][4] ) );
  OR2X1 U132 ( .A(\u_div/PartRem[51][2] ), .B(\u_div/PartRem[51][3] ), .Y(
        \u_div/u_add_PartRem_2_50/n3 ) );
  ADDHXL U133 ( .A(\u_div/PartRem[52][4] ), .B(\u_div/u_add_PartRem_2_51/n3 ), 
        .CO(\u_div/u_add_PartRem_2_51/n2 ), .S(\u_div/SumTmp[51][4] ) );
  OR2X1 U134 ( .A(\u_div/PartRem[52][2] ), .B(\u_div/PartRem[52][3] ), .Y(
        \u_div/u_add_PartRem_2_51/n3 ) );
  ADDHXL U135 ( .A(\u_div/PartRem[53][4] ), .B(\u_div/u_add_PartRem_2_52/n3 ), 
        .CO(\u_div/u_add_PartRem_2_52/n2 ), .S(\u_div/SumTmp[52][4] ) );
  ADDHXL U136 ( .A(\u_div/PartRem[54][4] ), .B(\u_div/u_add_PartRem_2_53/n3 ), 
        .CO(\u_div/u_add_PartRem_2_53/n2 ), .S(\u_div/SumTmp[53][4] ) );
  OR2X1 U137 ( .A(\u_div/PartRem[54][2] ), .B(\u_div/PartRem[54][3] ), .Y(
        \u_div/u_add_PartRem_2_53/n3 ) );
  ADDHXL U138 ( .A(\u_div/PartRem[55][4] ), .B(\u_div/u_add_PartRem_2_54/n3 ), 
        .CO(\u_div/u_add_PartRem_2_54/n2 ), .S(\u_div/SumTmp[54][4] ) );
  OR2X1 U139 ( .A(\u_div/PartRem[55][2] ), .B(\u_div/PartRem[55][3] ), .Y(
        \u_div/u_add_PartRem_2_54/n3 ) );
  ADDHXL U140 ( .A(\u_div/PartRem[56][4] ), .B(\u_div/u_add_PartRem_2_55/n3 ), 
        .CO(\u_div/u_add_PartRem_2_55/n2 ), .S(\u_div/SumTmp[55][4] ) );
  OR2X1 U141 ( .A(\u_div/PartRem[56][2] ), .B(\u_div/PartRem[56][3] ), .Y(
        \u_div/u_add_PartRem_2_55/n3 ) );
  ADDHXL U142 ( .A(\u_div/PartRem[57][4] ), .B(\u_div/u_add_PartRem_2_56/n3 ), 
        .CO(\u_div/u_add_PartRem_2_56/n2 ), .S(\u_div/SumTmp[56][4] ) );
  OR2X1 U143 ( .A(\u_div/PartRem[57][2] ), .B(\u_div/PartRem[57][3] ), .Y(
        \u_div/u_add_PartRem_2_56/n3 ) );
  ADDHXL U144 ( .A(\u_div/PartRem[58][4] ), .B(\u_div/u_add_PartRem_2_57/n3 ), 
        .CO(\u_div/u_add_PartRem_2_57/n2 ), .S(\u_div/SumTmp[57][4] ) );
  OR2X1 U145 ( .A(\u_div/PartRem[58][2] ), .B(\u_div/PartRem[58][3] ), .Y(
        \u_div/u_add_PartRem_2_57/n3 ) );
  OR2X1 U146 ( .A(\u_div/PartRem[59][2] ), .B(\u_div/PartRem[59][3] ), .Y(
        \u_div/u_add_PartRem_2_58/n3 ) );
  NOR2X1 U147 ( .A(\u_div/PartRem[63][0] ), .B(\u_div/PartRem[62][0] ), .Y(n8)
         );
  OR2X1 U148 ( .A(\u_div/PartRem[16][5] ), .B(\u_div/u_add_PartRem_2_15/n2 ), 
        .Y(\u_div/CryTmp[15][6] ) );
  OR2X1 U149 ( .A(\u_div/PartRem[21][5] ), .B(\u_div/u_add_PartRem_2_20/n2 ), 
        .Y(\u_div/CryTmp[20][6] ) );
  ADDHXL U150 ( .A(\u_div/PartRem[2][4] ), .B(\u_div/u_add_PartRem_2_1/n3 ), 
        .CO(\u_div/u_add_PartRem_2_1/n2 ), .S(\u_div/SumTmp[1][4] ) );
  OR2X1 U151 ( .A(\u_div/PartRem[2][2] ), .B(\u_div/PartRem[2][3] ), .Y(
        \u_div/u_add_PartRem_2_1/n3 ) );
  OR2X1 U152 ( .A(\u_div/PartRem[26][5] ), .B(\u_div/u_add_PartRem_2_25/n2 ), 
        .Y(\u_div/CryTmp[25][6] ) );
  OR2X1 U153 ( .A(\u_div/PartRem[31][5] ), .B(\u_div/u_add_PartRem_2_30/n2 ), 
        .Y(\u_div/CryTmp[30][6] ) );
  OR2X1 U154 ( .A(\u_div/PartRem[36][5] ), .B(\u_div/u_add_PartRem_2_35/n2 ), 
        .Y(\u_div/CryTmp[35][6] ) );
  OR2X1 U155 ( .A(\u_div/PartRem[41][5] ), .B(\u_div/u_add_PartRem_2_40/n2 ), 
        .Y(\u_div/CryTmp[40][6] ) );
  OR2X1 U156 ( .A(\u_div/PartRem[46][5] ), .B(\u_div/u_add_PartRem_2_45/n2 ), 
        .Y(\u_div/CryTmp[45][6] ) );
  OR2X1 U157 ( .A(\u_div/PartRem[51][5] ), .B(\u_div/u_add_PartRem_2_50/n2 ), 
        .Y(\u_div/CryTmp[50][6] ) );
  OR2X1 U158 ( .A(\u_div/PartRem[56][5] ), .B(\u_div/u_add_PartRem_2_55/n2 ), 
        .Y(\u_div/CryTmp[55][6] ) );
  NOR2BX2 U159 ( .AN(\u_div/PartRem[64][0] ), .B(n8), .Y(\u_div/CryTmp[59][6] ) );
  AO21X1 U160 ( .A0(\u_div/PartRem[1][4] ), .A1(n6), .B0(\u_div/PartRem[1][5] ), .Y(\u_div/CryTmp[0][6] ) );
  XNOR2XL U161 ( .A(\u_div/PartRem[64][0] ), .B(n8), .Y(\u_div/SumTmp[59][4] )
         );
  XOR2XL U162 ( .A(\u_div/CryTmp[59][6] ), .B(n3), .Y(\u_div/QInv[59] ) );
  XOR2XL U163 ( .A(\u_div/CryTmp[57][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[57] ) );
  XOR2XL U164 ( .A(\u_div/CryTmp[54][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[54] ) );
  XOR2XL U165 ( .A(\u_div/CryTmp[55][6] ), .B(n4), .Y(\u_div/QInv[55] ) );
  XOR2XL U166 ( .A(\u_div/CryTmp[52][6] ), .B(n4), .Y(\u_div/QInv[52] ) );
  XOR2XL U167 ( .A(\u_div/CryTmp[1][6] ), .B(n4), .Y(\u_div/QInv[1] ) );
  XOR2XL U168 ( .A(\u_div/CryTmp[51][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[51] ) );
  XOR2XL U169 ( .A(\u_div/CryTmp[46][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[46] ) );
  XOR2XL U170 ( .A(\u_div/CryTmp[43][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[43] ) );
  XOR2XL U171 ( .A(\u_div/CryTmp[47][6] ), .B(n4), .Y(\u_div/QInv[47] ) );
  XOR2XL U172 ( .A(\u_div/CryTmp[44][6] ), .B(n4), .Y(\u_div/QInv[44] ) );
  XOR2XL U173 ( .A(\u_div/CryTmp[40][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[40] ) );
  XOR2XL U174 ( .A(\u_div/CryTmp[41][6] ), .B(n4), .Y(\u_div/QInv[41] ) );
  XOR2XL U175 ( .A(\u_div/CryTmp[35][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[35] ) );
  XOR2XL U176 ( .A(\u_div/CryTmp[34][6] ), .B(n4), .Y(\u_div/QInv[34] ) );
  XOR2XL U177 ( .A(\u_div/CryTmp[36][6] ), .B(n4), .Y(\u_div/QInv[36] ) );
  XOR2XL U178 ( .A(\u_div/CryTmp[33][6] ), .B(n5), .Y(\u_div/QInv[33] ) );
  XOR2XL U179 ( .A(\u_div/CryTmp[30][6] ), .B(n5), .Y(\u_div/QInv[30] ) );
  XOR2XL U180 ( .A(\u_div/CryTmp[31][6] ), .B(n4), .Y(\u_div/QInv[31] ) );
  XOR2XL U181 ( .A(\u_div/CryTmp[25][6] ), .B(n5), .Y(\u_div/QInv[25] ) );
  XOR2XL U182 ( .A(\u_div/CryTmp[26][6] ), .B(n4), .Y(\u_div/QInv[26] ) );
  XOR2XL U183 ( .A(\u_div/CryTmp[23][6] ), .B(n4), .Y(\u_div/QInv[23] ) );
  XOR2XL U184 ( .A(\u_div/CryTmp[22][6] ), .B(n5), .Y(\u_div/QInv[22] ) );
  XOR2XL U185 ( .A(\u_div/CryTmp[20][6] ), .B(n4), .Y(\u_div/QInv[20] ) );
  XOR2XL U186 ( .A(\u_div/CryTmp[17][6] ), .B(n5), .Y(\u_div/QInv[17] ) );
  XOR2XL U187 ( .A(\u_div/CryTmp[16][6] ), .B(n4), .Y(\u_div/QInv[16] ) );
  XOR2XL U188 ( .A(\u_div/CryTmp[15][6] ), .B(n3), .Y(\u_div/QInv[15] ) );
  XOR2XL U189 ( .A(\u_div/CryTmp[14][6] ), .B(n4), .Y(\u_div/QInv[14] ) );
  XOR2XL U190 ( .A(\u_div/CryTmp[11][6] ), .B(n4), .Y(\u_div/QInv[11] ) );
  XOR2XL U191 ( .A(\u_div/CryTmp[12][6] ), .B(n4), .Y(\u_div/QInv[12] ) );
  XOR2XL U192 ( .A(\u_div/CryTmp[4][6] ), .B(n4), .Y(\u_div/QInv[4] ) );
  XOR2XL U193 ( .A(\u_div/CryTmp[5][6] ), .B(n4), .Y(\u_div/QInv[5] ) );
  XOR2XL U194 ( .A(\u_div/CryTmp[6][6] ), .B(n4), .Y(\u_div/QInv[6] ) );
  XOR2XL U195 ( .A(\u_div/CryTmp[7][6] ), .B(n4), .Y(\u_div/QInv[7] ) );
  XOR2XL U196 ( .A(\u_div/CryTmp[10][6] ), .B(n4), .Y(\u_div/QInv[10] ) );
  XOR2XL U197 ( .A(\u_div/CryTmp[13][6] ), .B(n4), .Y(\u_div/QInv[13] ) );
  XOR2XL U198 ( .A(\u_div/CryTmp[53][6] ), .B(n3), .Y(\u_div/QInv[53] ) );
  XOR2XL U199 ( .A(\u_div/CryTmp[50][6] ), .B(n3), .Y(\u_div/QInv[50] ) );
  XOR2XL U200 ( .A(\u_div/CryTmp[45][6] ), .B(n3), .Y(\u_div/QInv[45] ) );
  XOR2XL U201 ( .A(\u_div/CryTmp[42][6] ), .B(n3), .Y(\u_div/QInv[42] ) );
  XOR2XL U202 ( .A(\u_div/CryTmp[37][6] ), .B(n3), .Y(\u_div/QInv[37] ) );
  XOR2XL U203 ( .A(\u_div/CryTmp[32][6] ), .B(n3), .Y(\u_div/QInv[32] ) );
  XOR2XL U204 ( .A(\u_div/CryTmp[27][6] ), .B(n3), .Y(\u_div/QInv[27] ) );
  XOR2XL U205 ( .A(\u_div/CryTmp[24][6] ), .B(n3), .Y(\u_div/QInv[24] ) );
  XOR2XL U206 ( .A(\u_div/CryTmp[21][6] ), .B(n3), .Y(\u_div/QInv[21] ) );
  XOR2XL U207 ( .A(\u_div/CryTmp[2][6] ), .B(n3), .Y(\u_div/QInv[2] ) );
  XOR2XL U208 ( .A(\u_div/CryTmp[3][6] ), .B(n3), .Y(\u_div/QInv[3] ) );
  INVXL U209 ( .A(\u_div/PartRem[59][2] ), .Y(\u_div/SumTmp[58][2] ) );
  INVXL U210 ( .A(\u_div/PartRem[55][2] ), .Y(\u_div/SumTmp[54][2] ) );
  INVXL U211 ( .A(\u_div/PartRem[50][2] ), .Y(\u_div/SumTmp[49][2] ) );
  INVXL U212 ( .A(\u_div/PartRem[45][2] ), .Y(\u_div/SumTmp[44][2] ) );
  INVXL U213 ( .A(\u_div/PartRem[40][2] ), .Y(\u_div/SumTmp[39][2] ) );
  INVXL U214 ( .A(\u_div/PartRem[35][2] ), .Y(\u_div/SumTmp[34][2] ) );
  INVXL U215 ( .A(\u_div/PartRem[30][2] ), .Y(\u_div/SumTmp[29][2] ) );
  INVXL U216 ( .A(\u_div/PartRem[25][2] ), .Y(\u_div/SumTmp[24][2] ) );
  INVXL U217 ( .A(\u_div/PartRem[20][2] ), .Y(\u_div/SumTmp[19][2] ) );
  INVXL U218 ( .A(\u_div/PartRem[15][2] ), .Y(\u_div/SumTmp[14][2] ) );
  INVXL U219 ( .A(\u_div/PartRem[10][2] ), .Y(\u_div/SumTmp[9][2] ) );
  INVXL U220 ( .A(\u_div/PartRem[5][2] ), .Y(\u_div/SumTmp[4][2] ) );
  INVX3 U221 ( .A(n2), .Y(n3) );
  MXI2X1 U222 ( .A(\u_div/SumTmp[1][1] ), .B(\u_div/SumTmp[1][1] ), .S0(
        \u_div/CryTmp[1][6] ), .Y(n1) );
  CLKINVX1 U223 ( .A(n5), .Y(n2) );
  MXI2X1 U224 ( .A(n7), .B(\u_div/PartRem[62][0] ), .S0(\u_div/CryTmp[59][6] ), 
        .Y(\u_div/PartRem[59][3] ) );
  CLKINVX1 U225 ( .A(\u_div/PartRem[62][0] ), .Y(n7) );
  MXI2X1 U226 ( .A(\u_div/SumTmp[58][2] ), .B(\u_div/PartRem[59][2] ), .S0(
        \u_div/CryTmp[58][6] ), .Y(\u_div/PartRem[58][3] ) );
  MXI2X1 U227 ( .A(\u_div/SumTmp[57][2] ), .B(\u_div/PartRem[58][2] ), .S0(
        \u_div/CryTmp[57][6] ), .Y(\u_div/PartRem[57][3] ) );
  CLKINVX1 U228 ( .A(\u_div/PartRem[58][2] ), .Y(\u_div/SumTmp[57][2] ) );
  CLKINVX1 U229 ( .A(\u_div/PartRem[57][2] ), .Y(\u_div/SumTmp[56][2] ) );
  MXI2X1 U230 ( .A(\u_div/SumTmp[54][2] ), .B(\u_div/PartRem[55][2] ), .S0(
        \u_div/CryTmp[54][6] ), .Y(\u_div/PartRem[54][3] ) );
  CLKINVX1 U231 ( .A(\u_div/PartRem[54][2] ), .Y(\u_div/SumTmp[53][2] ) );
  MXI2X1 U232 ( .A(\u_div/SumTmp[52][2] ), .B(\u_div/PartRem[53][2] ), .S0(
        \u_div/CryTmp[52][6] ), .Y(\u_div/PartRem[52][3] ) );
  CLKINVX1 U233 ( .A(\u_div/PartRem[53][2] ), .Y(\u_div/SumTmp[52][2] ) );
  MXI2X1 U234 ( .A(\u_div/SumTmp[51][2] ), .B(\u_div/PartRem[52][2] ), .S0(
        \u_div/CryTmp[51][6] ), .Y(\u_div/PartRem[51][3] ) );
  CLKINVX1 U235 ( .A(\u_div/PartRem[52][2] ), .Y(\u_div/SumTmp[51][2] ) );
  CLKINVX1 U236 ( .A(\u_div/PartRem[49][2] ), .Y(\u_div/SumTmp[48][2] ) );
  MXI2X1 U237 ( .A(\u_div/SumTmp[47][2] ), .B(\u_div/PartRem[48][2] ), .S0(
        \u_div/CryTmp[47][6] ), .Y(\u_div/PartRem[47][3] ) );
  CLKINVX1 U238 ( .A(\u_div/PartRem[48][2] ), .Y(\u_div/SumTmp[47][2] ) );
  MXI2X1 U239 ( .A(\u_div/SumTmp[46][2] ), .B(\u_div/PartRem[47][2] ), .S0(
        \u_div/CryTmp[46][6] ), .Y(\u_div/PartRem[46][3] ) );
  CLKINVX1 U240 ( .A(\u_div/PartRem[47][2] ), .Y(\u_div/SumTmp[46][2] ) );
  MXI2X1 U241 ( .A(\u_div/SumTmp[44][2] ), .B(\u_div/PartRem[45][2] ), .S0(
        \u_div/CryTmp[44][6] ), .Y(\u_div/PartRem[44][3] ) );
  CLKINVX1 U242 ( .A(\u_div/PartRem[44][2] ), .Y(\u_div/SumTmp[43][2] ) );
  MXI2X1 U243 ( .A(\u_div/SumTmp[42][2] ), .B(\u_div/PartRem[43][2] ), .S0(
        \u_div/CryTmp[42][6] ), .Y(\u_div/PartRem[42][3] ) );
  CLKINVX1 U244 ( .A(\u_div/PartRem[43][2] ), .Y(\u_div/SumTmp[42][2] ) );
  MXI2X1 U245 ( .A(\u_div/SumTmp[41][2] ), .B(\u_div/PartRem[42][2] ), .S0(
        \u_div/CryTmp[41][6] ), .Y(\u_div/PartRem[41][3] ) );
  CLKINVX1 U246 ( .A(\u_div/PartRem[42][2] ), .Y(\u_div/SumTmp[41][2] ) );
  MXI2X1 U247 ( .A(\u_div/SumTmp[39][2] ), .B(\u_div/PartRem[40][2] ), .S0(
        \u_div/CryTmp[39][6] ), .Y(\u_div/PartRem[39][3] ) );
  CLKINVX1 U248 ( .A(\u_div/PartRem[39][2] ), .Y(\u_div/SumTmp[38][2] ) );
  MXI2X1 U249 ( .A(\u_div/SumTmp[37][2] ), .B(\u_div/PartRem[38][2] ), .S0(
        \u_div/CryTmp[37][6] ), .Y(\u_div/PartRem[37][3] ) );
  CLKINVX1 U250 ( .A(\u_div/PartRem[38][2] ), .Y(\u_div/SumTmp[37][2] ) );
  MXI2X1 U251 ( .A(\u_div/SumTmp[36][2] ), .B(\u_div/PartRem[37][2] ), .S0(
        \u_div/CryTmp[36][6] ), .Y(\u_div/PartRem[36][3] ) );
  CLKINVX1 U252 ( .A(\u_div/PartRem[37][2] ), .Y(\u_div/SumTmp[36][2] ) );
  MXI2X1 U253 ( .A(\u_div/SumTmp[34][2] ), .B(\u_div/PartRem[35][2] ), .S0(
        \u_div/CryTmp[34][6] ), .Y(\u_div/PartRem[34][3] ) );
  CLKINVX1 U254 ( .A(\u_div/PartRem[34][2] ), .Y(\u_div/SumTmp[33][2] ) );
  MXI2X1 U255 ( .A(\u_div/SumTmp[32][2] ), .B(\u_div/PartRem[33][2] ), .S0(
        \u_div/CryTmp[32][6] ), .Y(\u_div/PartRem[32][3] ) );
  CLKINVX1 U256 ( .A(\u_div/PartRem[33][2] ), .Y(\u_div/SumTmp[32][2] ) );
  MXI2X1 U257 ( .A(\u_div/SumTmp[31][2] ), .B(\u_div/PartRem[32][2] ), .S0(
        \u_div/CryTmp[31][6] ), .Y(\u_div/PartRem[31][3] ) );
  CLKINVX1 U258 ( .A(\u_div/PartRem[32][2] ), .Y(\u_div/SumTmp[31][2] ) );
  MXI2X1 U259 ( .A(\u_div/SumTmp[29][2] ), .B(\u_div/PartRem[30][2] ), .S0(
        \u_div/CryTmp[29][6] ), .Y(\u_div/PartRem[29][3] ) );
  CLKINVX1 U260 ( .A(\u_div/PartRem[29][2] ), .Y(\u_div/SumTmp[28][2] ) );
  MXI2X1 U261 ( .A(\u_div/SumTmp[27][2] ), .B(\u_div/PartRem[28][2] ), .S0(
        \u_div/CryTmp[27][6] ), .Y(\u_div/PartRem[27][3] ) );
  CLKINVX1 U262 ( .A(\u_div/PartRem[28][2] ), .Y(\u_div/SumTmp[27][2] ) );
  MXI2X1 U263 ( .A(\u_div/SumTmp[26][2] ), .B(\u_div/PartRem[27][2] ), .S0(
        \u_div/CryTmp[26][6] ), .Y(\u_div/PartRem[26][3] ) );
  CLKINVX1 U264 ( .A(\u_div/PartRem[27][2] ), .Y(\u_div/SumTmp[26][2] ) );
  MXI2X1 U265 ( .A(\u_div/SumTmp[24][2] ), .B(\u_div/PartRem[25][2] ), .S0(
        \u_div/CryTmp[24][6] ), .Y(\u_div/PartRem[24][3] ) );
  CLKINVX1 U266 ( .A(\u_div/PartRem[24][2] ), .Y(\u_div/SumTmp[23][2] ) );
  MXI2X1 U267 ( .A(\u_div/SumTmp[22][2] ), .B(\u_div/PartRem[23][2] ), .S0(
        \u_div/CryTmp[22][6] ), .Y(\u_div/PartRem[22][3] ) );
  CLKINVX1 U268 ( .A(\u_div/PartRem[23][2] ), .Y(\u_div/SumTmp[22][2] ) );
  MXI2X1 U269 ( .A(\u_div/SumTmp[21][2] ), .B(\u_div/PartRem[22][2] ), .S0(
        \u_div/CryTmp[21][6] ), .Y(\u_div/PartRem[21][3] ) );
  CLKINVX1 U270 ( .A(\u_div/PartRem[22][2] ), .Y(\u_div/SumTmp[21][2] ) );
  CLKINVX1 U271 ( .A(\u_div/PartRem[19][2] ), .Y(\u_div/SumTmp[18][2] ) );
  MXI2X1 U272 ( .A(\u_div/SumTmp[17][2] ), .B(\u_div/PartRem[18][2] ), .S0(
        \u_div/CryTmp[17][6] ), .Y(\u_div/PartRem[17][3] ) );
  CLKINVX1 U273 ( .A(\u_div/PartRem[18][2] ), .Y(\u_div/SumTmp[17][2] ) );
  MXI2X1 U274 ( .A(\u_div/SumTmp[16][2] ), .B(\u_div/PartRem[17][2] ), .S0(
        \u_div/CryTmp[16][6] ), .Y(\u_div/PartRem[16][3] ) );
  CLKINVX1 U275 ( .A(\u_div/PartRem[17][2] ), .Y(\u_div/SumTmp[16][2] ) );
  MXI2X1 U276 ( .A(\u_div/SumTmp[14][2] ), .B(\u_div/PartRem[15][2] ), .S0(
        \u_div/CryTmp[14][6] ), .Y(\u_div/PartRem[14][3] ) );
  CLKINVX1 U277 ( .A(\u_div/PartRem[14][2] ), .Y(\u_div/SumTmp[13][2] ) );
  MXI2X1 U278 ( .A(\u_div/SumTmp[12][2] ), .B(\u_div/PartRem[13][2] ), .S0(
        \u_div/CryTmp[12][6] ), .Y(\u_div/PartRem[12][3] ) );
  CLKINVX1 U279 ( .A(\u_div/PartRem[13][2] ), .Y(\u_div/SumTmp[12][2] ) );
  MXI2X1 U280 ( .A(\u_div/SumTmp[11][2] ), .B(\u_div/PartRem[12][2] ), .S0(
        \u_div/CryTmp[11][6] ), .Y(\u_div/PartRem[11][3] ) );
  CLKINVX1 U281 ( .A(\u_div/PartRem[12][2] ), .Y(\u_div/SumTmp[11][2] ) );
  CLKINVX1 U282 ( .A(\u_div/PartRem[9][2] ), .Y(\u_div/SumTmp[8][2] ) );
  CLKINVX1 U283 ( .A(\u_div/PartRem[8][2] ), .Y(\u_div/SumTmp[7][2] ) );
  MXI2X1 U284 ( .A(\u_div/SumTmp[6][2] ), .B(\u_div/PartRem[7][2] ), .S0(
        \u_div/CryTmp[6][6] ), .Y(\u_div/PartRem[6][3] ) );
  CLKINVX1 U285 ( .A(\u_div/PartRem[7][2] ), .Y(\u_div/SumTmp[6][2] ) );
  MXI2X1 U286 ( .A(\u_div/SumTmp[4][2] ), .B(\u_div/PartRem[5][2] ), .S0(
        \u_div/CryTmp[4][6] ), .Y(\u_div/PartRem[4][3] ) );
  CLKINVX1 U287 ( .A(\u_div/PartRem[4][2] ), .Y(\u_div/SumTmp[3][2] ) );
  MXI2X1 U288 ( .A(\u_div/SumTmp[2][2] ), .B(\u_div/PartRem[3][2] ), .S0(
        \u_div/CryTmp[2][6] ), .Y(\u_div/PartRem[2][3] ) );
  CLKINVX1 U289 ( .A(\u_div/PartRem[3][2] ), .Y(\u_div/SumTmp[2][2] ) );
  MXI2X1 U290 ( .A(\u_div/SumTmp[55][2] ), .B(\u_div/PartRem[56][2] ), .S0(
        \u_div/CryTmp[55][6] ), .Y(\u_div/PartRem[55][3] ) );
  CLKINVX1 U291 ( .A(\u_div/PartRem[56][2] ), .Y(\u_div/SumTmp[55][2] ) );
  MXI2X1 U292 ( .A(\u_div/SumTmp[50][2] ), .B(\u_div/PartRem[51][2] ), .S0(
        \u_div/CryTmp[50][6] ), .Y(\u_div/PartRem[50][3] ) );
  CLKINVX1 U293 ( .A(\u_div/PartRem[51][2] ), .Y(\u_div/SumTmp[50][2] ) );
  MXI2X1 U294 ( .A(\u_div/SumTmp[45][2] ), .B(\u_div/PartRem[46][2] ), .S0(
        \u_div/CryTmp[45][6] ), .Y(\u_div/PartRem[45][3] ) );
  CLKINVX1 U295 ( .A(\u_div/PartRem[46][2] ), .Y(\u_div/SumTmp[45][2] ) );
  MXI2X1 U296 ( .A(\u_div/SumTmp[40][2] ), .B(\u_div/PartRem[41][2] ), .S0(
        \u_div/CryTmp[40][6] ), .Y(\u_div/PartRem[40][3] ) );
  CLKINVX1 U297 ( .A(\u_div/PartRem[41][2] ), .Y(\u_div/SumTmp[40][2] ) );
  MXI2X1 U298 ( .A(\u_div/SumTmp[35][2] ), .B(\u_div/PartRem[36][2] ), .S0(
        \u_div/CryTmp[35][6] ), .Y(\u_div/PartRem[35][3] ) );
  CLKINVX1 U299 ( .A(\u_div/PartRem[36][2] ), .Y(\u_div/SumTmp[35][2] ) );
  MXI2X1 U300 ( .A(\u_div/SumTmp[30][2] ), .B(\u_div/PartRem[31][2] ), .S0(
        \u_div/CryTmp[30][6] ), .Y(\u_div/PartRem[30][3] ) );
  CLKINVX1 U301 ( .A(\u_div/PartRem[31][2] ), .Y(\u_div/SumTmp[30][2] ) );
  MXI2X1 U302 ( .A(\u_div/SumTmp[25][2] ), .B(\u_div/PartRem[26][2] ), .S0(
        \u_div/CryTmp[25][6] ), .Y(\u_div/PartRem[25][3] ) );
  CLKINVX1 U303 ( .A(\u_div/PartRem[26][2] ), .Y(\u_div/SumTmp[25][2] ) );
  MXI2X1 U304 ( .A(\u_div/SumTmp[20][2] ), .B(\u_div/PartRem[21][2] ), .S0(
        \u_div/CryTmp[20][6] ), .Y(\u_div/PartRem[20][3] ) );
  CLKINVX1 U305 ( .A(\u_div/PartRem[21][2] ), .Y(\u_div/SumTmp[20][2] ) );
  MXI2X1 U306 ( .A(\u_div/SumTmp[15][2] ), .B(\u_div/PartRem[16][2] ), .S0(
        \u_div/CryTmp[15][6] ), .Y(\u_div/PartRem[15][3] ) );
  CLKINVX1 U307 ( .A(\u_div/PartRem[16][2] ), .Y(\u_div/SumTmp[15][2] ) );
  MXI2X1 U308 ( .A(\u_div/SumTmp[10][2] ), .B(\u_div/PartRem[11][2] ), .S0(
        \u_div/CryTmp[10][6] ), .Y(\u_div/PartRem[10][3] ) );
  CLKINVX1 U309 ( .A(\u_div/PartRem[11][2] ), .Y(\u_div/SumTmp[10][2] ) );
  MXI2X1 U310 ( .A(\u_div/SumTmp[5][2] ), .B(\u_div/PartRem[6][2] ), .S0(
        \u_div/CryTmp[5][6] ), .Y(\u_div/PartRem[5][3] ) );
  CLKINVX1 U311 ( .A(\u_div/PartRem[6][2] ), .Y(\u_div/SumTmp[5][2] ) );
  CLKINVX1 U312 ( .A(\u_div/PartRem[2][2] ), .Y(\u_div/SumTmp[1][2] ) );
  INVX4 U313 ( .A(n2), .Y(n4) );
  CLKBUFX3 U314 ( .A(\u_div/QInv[63] ), .Y(n5) );
  XNOR2X1 U315 ( .A(\u_div/PartRem[59][3] ), .B(\u_div/PartRem[59][2] ), .Y(
        \u_div/SumTmp[58][3] ) );
  OR2X1 U316 ( .A(\u_div/PartRem[58][5] ), .B(\u_div/u_add_PartRem_2_57/n2 ), 
        .Y(\u_div/CryTmp[57][6] ) );
  XNOR2X1 U317 ( .A(\u_div/PartRem[58][3] ), .B(\u_div/PartRem[58][2] ), .Y(
        \u_div/SumTmp[57][3] ) );
  XNOR2X1 U318 ( .A(\u_div/PartRem[57][3] ), .B(\u_div/PartRem[57][2] ), .Y(
        \u_div/SumTmp[56][3] ) );
  XNOR2X1 U319 ( .A(\u_div/PartRem[56][3] ), .B(\u_div/PartRem[56][2] ), .Y(
        \u_div/SumTmp[55][3] ) );
  OR2X1 U320 ( .A(\u_div/PartRem[55][5] ), .B(\u_div/u_add_PartRem_2_54/n2 ), 
        .Y(\u_div/CryTmp[54][6] ) );
  XNOR2X1 U321 ( .A(\u_div/PartRem[55][3] ), .B(\u_div/PartRem[55][2] ), .Y(
        \u_div/SumTmp[54][3] ) );
  OR2X1 U322 ( .A(\u_div/PartRem[54][5] ), .B(\u_div/u_add_PartRem_2_53/n2 ), 
        .Y(\u_div/CryTmp[53][6] ) );
  XNOR2X1 U323 ( .A(\u_div/PartRem[54][3] ), .B(\u_div/PartRem[54][2] ), .Y(
        \u_div/SumTmp[53][3] ) );
  OR2X1 U324 ( .A(\u_div/PartRem[53][5] ), .B(\u_div/u_add_PartRem_2_52/n2 ), 
        .Y(\u_div/CryTmp[52][6] ) );
  XNOR2X1 U325 ( .A(\u_div/PartRem[53][3] ), .B(\u_div/PartRem[53][2] ), .Y(
        \u_div/SumTmp[52][3] ) );
  OR2X1 U326 ( .A(\u_div/PartRem[53][2] ), .B(\u_div/PartRem[53][3] ), .Y(
        \u_div/u_add_PartRem_2_52/n3 ) );
  OR2X1 U327 ( .A(\u_div/PartRem[52][5] ), .B(\u_div/u_add_PartRem_2_51/n2 ), 
        .Y(\u_div/CryTmp[51][6] ) );
  XNOR2X1 U328 ( .A(\u_div/PartRem[52][3] ), .B(\u_div/PartRem[52][2] ), .Y(
        \u_div/SumTmp[51][3] ) );
  XNOR2X1 U329 ( .A(\u_div/PartRem[51][3] ), .B(\u_div/PartRem[51][2] ), .Y(
        \u_div/SumTmp[50][3] ) );
  XNOR2X1 U330 ( .A(\u_div/PartRem[50][3] ), .B(\u_div/PartRem[50][2] ), .Y(
        \u_div/SumTmp[49][3] ) );
  XNOR2X1 U331 ( .A(\u_div/PartRem[49][3] ), .B(\u_div/PartRem[49][2] ), .Y(
        \u_div/SumTmp[48][3] ) );
  OR2X1 U332 ( .A(\u_div/PartRem[48][5] ), .B(\u_div/u_add_PartRem_2_47/n2 ), 
        .Y(\u_div/CryTmp[47][6] ) );
  XNOR2X1 U333 ( .A(\u_div/PartRem[48][3] ), .B(\u_div/PartRem[48][2] ), .Y(
        \u_div/SumTmp[47][3] ) );
  OR2X1 U334 ( .A(\u_div/PartRem[48][2] ), .B(\u_div/PartRem[48][3] ), .Y(
        \u_div/u_add_PartRem_2_47/n3 ) );
  OR2X1 U335 ( .A(\u_div/PartRem[47][5] ), .B(\u_div/u_add_PartRem_2_46/n2 ), 
        .Y(\u_div/CryTmp[46][6] ) );
  XNOR2X1 U336 ( .A(\u_div/PartRem[47][3] ), .B(\u_div/PartRem[47][2] ), .Y(
        \u_div/SumTmp[46][3] ) );
  XNOR2X1 U337 ( .A(\u_div/PartRem[46][3] ), .B(\u_div/PartRem[46][2] ), .Y(
        \u_div/SumTmp[45][3] ) );
  OR2X1 U338 ( .A(\u_div/PartRem[45][5] ), .B(\u_div/u_add_PartRem_2_44/n2 ), 
        .Y(\u_div/CryTmp[44][6] ) );
  XNOR2X1 U339 ( .A(\u_div/PartRem[45][3] ), .B(\u_div/PartRem[45][2] ), .Y(
        \u_div/SumTmp[44][3] ) );
  OR2X1 U340 ( .A(\u_div/PartRem[44][5] ), .B(\u_div/u_add_PartRem_2_43/n2 ), 
        .Y(\u_div/CryTmp[43][6] ) );
  XNOR2X1 U341 ( .A(\u_div/PartRem[44][3] ), .B(\u_div/PartRem[44][2] ), .Y(
        \u_div/SumTmp[43][3] ) );
  OR2X1 U342 ( .A(\u_div/PartRem[43][5] ), .B(\u_div/u_add_PartRem_2_42/n2 ), 
        .Y(\u_div/CryTmp[42][6] ) );
  XNOR2X1 U343 ( .A(\u_div/PartRem[43][3] ), .B(\u_div/PartRem[43][2] ), .Y(
        \u_div/SumTmp[42][3] ) );
  OR2X1 U344 ( .A(\u_div/PartRem[43][2] ), .B(\u_div/PartRem[43][3] ), .Y(
        \u_div/u_add_PartRem_2_42/n3 ) );
  OR2X1 U345 ( .A(\u_div/PartRem[42][5] ), .B(\u_div/u_add_PartRem_2_41/n2 ), 
        .Y(\u_div/CryTmp[41][6] ) );
  XNOR2X1 U346 ( .A(\u_div/PartRem[42][3] ), .B(\u_div/PartRem[42][2] ), .Y(
        \u_div/SumTmp[41][3] ) );
  XNOR2X1 U347 ( .A(\u_div/PartRem[41][3] ), .B(\u_div/PartRem[41][2] ), .Y(
        \u_div/SumTmp[40][3] ) );
  XNOR2X1 U348 ( .A(\u_div/PartRem[40][3] ), .B(\u_div/PartRem[40][2] ), .Y(
        \u_div/SumTmp[39][3] ) );
  XNOR2X1 U349 ( .A(\u_div/PartRem[39][3] ), .B(\u_div/PartRem[39][2] ), .Y(
        \u_div/SumTmp[38][3] ) );
  OR2X1 U350 ( .A(\u_div/PartRem[38][5] ), .B(\u_div/u_add_PartRem_2_37/n2 ), 
        .Y(\u_div/CryTmp[37][6] ) );
  XNOR2X1 U351 ( .A(\u_div/PartRem[38][3] ), .B(\u_div/PartRem[38][2] ), .Y(
        \u_div/SumTmp[37][3] ) );
  OR2X1 U352 ( .A(\u_div/PartRem[38][2] ), .B(\u_div/PartRem[38][3] ), .Y(
        \u_div/u_add_PartRem_2_37/n3 ) );
  OR2X1 U353 ( .A(\u_div/PartRem[37][5] ), .B(\u_div/u_add_PartRem_2_36/n2 ), 
        .Y(\u_div/CryTmp[36][6] ) );
  XNOR2X1 U354 ( .A(\u_div/PartRem[37][3] ), .B(\u_div/PartRem[37][2] ), .Y(
        \u_div/SumTmp[36][3] ) );
  XNOR2X1 U355 ( .A(\u_div/PartRem[36][3] ), .B(\u_div/PartRem[36][2] ), .Y(
        \u_div/SumTmp[35][3] ) );
  OR2X1 U356 ( .A(\u_div/PartRem[35][5] ), .B(\u_div/u_add_PartRem_2_34/n2 ), 
        .Y(\u_div/CryTmp[34][6] ) );
  XNOR2X1 U357 ( .A(\u_div/PartRem[35][3] ), .B(\u_div/PartRem[35][2] ), .Y(
        \u_div/SumTmp[34][3] ) );
  OR2X1 U358 ( .A(\u_div/PartRem[34][5] ), .B(\u_div/u_add_PartRem_2_33/n2 ), 
        .Y(\u_div/CryTmp[33][6] ) );
  XNOR2X1 U359 ( .A(\u_div/PartRem[34][3] ), .B(\u_div/PartRem[34][2] ), .Y(
        \u_div/SumTmp[33][3] ) );
  OR2X1 U360 ( .A(\u_div/PartRem[33][5] ), .B(\u_div/u_add_PartRem_2_32/n2 ), 
        .Y(\u_div/CryTmp[32][6] ) );
  XNOR2X1 U361 ( .A(\u_div/PartRem[33][3] ), .B(\u_div/PartRem[33][2] ), .Y(
        \u_div/SumTmp[32][3] ) );
  OR2X1 U362 ( .A(\u_div/PartRem[33][2] ), .B(\u_div/PartRem[33][3] ), .Y(
        \u_div/u_add_PartRem_2_32/n3 ) );
  OR2X1 U363 ( .A(\u_div/PartRem[32][5] ), .B(\u_div/u_add_PartRem_2_31/n2 ), 
        .Y(\u_div/CryTmp[31][6] ) );
  XNOR2X1 U364 ( .A(\u_div/PartRem[32][3] ), .B(\u_div/PartRem[32][2] ), .Y(
        \u_div/SumTmp[31][3] ) );
  XNOR2X1 U365 ( .A(\u_div/PartRem[31][3] ), .B(\u_div/PartRem[31][2] ), .Y(
        \u_div/SumTmp[30][3] ) );
  XNOR2X1 U366 ( .A(\u_div/PartRem[30][3] ), .B(\u_div/PartRem[30][2] ), .Y(
        \u_div/SumTmp[29][3] ) );
  XNOR2X1 U367 ( .A(\u_div/PartRem[29][3] ), .B(\u_div/PartRem[29][2] ), .Y(
        \u_div/SumTmp[28][3] ) );
  OR2X1 U368 ( .A(\u_div/PartRem[28][5] ), .B(\u_div/u_add_PartRem_2_27/n2 ), 
        .Y(\u_div/CryTmp[27][6] ) );
  XNOR2X1 U369 ( .A(\u_div/PartRem[28][3] ), .B(\u_div/PartRem[28][2] ), .Y(
        \u_div/SumTmp[27][3] ) );
  OR2X1 U370 ( .A(\u_div/PartRem[28][2] ), .B(\u_div/PartRem[28][3] ), .Y(
        \u_div/u_add_PartRem_2_27/n3 ) );
  OR2X1 U371 ( .A(\u_div/PartRem[27][5] ), .B(\u_div/u_add_PartRem_2_26/n2 ), 
        .Y(\u_div/CryTmp[26][6] ) );
  XNOR2X1 U372 ( .A(\u_div/PartRem[27][3] ), .B(\u_div/PartRem[27][2] ), .Y(
        \u_div/SumTmp[26][3] ) );
  XNOR2X1 U373 ( .A(\u_div/PartRem[26][3] ), .B(\u_div/PartRem[26][2] ), .Y(
        \u_div/SumTmp[25][3] ) );
  OR2X1 U374 ( .A(\u_div/PartRem[25][5] ), .B(\u_div/u_add_PartRem_2_24/n2 ), 
        .Y(\u_div/CryTmp[24][6] ) );
  XNOR2X1 U375 ( .A(\u_div/PartRem[25][3] ), .B(\u_div/PartRem[25][2] ), .Y(
        \u_div/SumTmp[24][3] ) );
  OR2X1 U376 ( .A(\u_div/PartRem[24][5] ), .B(\u_div/u_add_PartRem_2_23/n2 ), 
        .Y(\u_div/CryTmp[23][6] ) );
  XNOR2X1 U377 ( .A(\u_div/PartRem[24][3] ), .B(\u_div/PartRem[24][2] ), .Y(
        \u_div/SumTmp[23][3] ) );
  OR2X1 U378 ( .A(\u_div/PartRem[23][5] ), .B(\u_div/u_add_PartRem_2_22/n2 ), 
        .Y(\u_div/CryTmp[22][6] ) );
  XNOR2X1 U379 ( .A(\u_div/PartRem[23][3] ), .B(\u_div/PartRem[23][2] ), .Y(
        \u_div/SumTmp[22][3] ) );
  OR2X1 U380 ( .A(\u_div/PartRem[23][2] ), .B(\u_div/PartRem[23][3] ), .Y(
        \u_div/u_add_PartRem_2_22/n3 ) );
  OR2X1 U381 ( .A(\u_div/PartRem[22][5] ), .B(\u_div/u_add_PartRem_2_21/n2 ), 
        .Y(\u_div/CryTmp[21][6] ) );
  XNOR2X1 U382 ( .A(\u_div/PartRem[22][3] ), .B(\u_div/PartRem[22][2] ), .Y(
        \u_div/SumTmp[21][3] ) );
  XNOR2X1 U383 ( .A(\u_div/PartRem[21][3] ), .B(\u_div/PartRem[21][2] ), .Y(
        \u_div/SumTmp[20][3] ) );
  XNOR2X1 U384 ( .A(\u_div/PartRem[20][3] ), .B(\u_div/PartRem[20][2] ), .Y(
        \u_div/SumTmp[19][3] ) );
  XNOR2X1 U385 ( .A(\u_div/PartRem[19][3] ), .B(\u_div/PartRem[19][2] ), .Y(
        \u_div/SumTmp[18][3] ) );
  OR2X1 U386 ( .A(\u_div/PartRem[18][5] ), .B(\u_div/u_add_PartRem_2_17/n2 ), 
        .Y(\u_div/CryTmp[17][6] ) );
  XNOR2X1 U387 ( .A(\u_div/PartRem[18][3] ), .B(\u_div/PartRem[18][2] ), .Y(
        \u_div/SumTmp[17][3] ) );
  OR2X1 U388 ( .A(\u_div/PartRem[18][2] ), .B(\u_div/PartRem[18][3] ), .Y(
        \u_div/u_add_PartRem_2_17/n3 ) );
  OR2X1 U389 ( .A(\u_div/PartRem[17][5] ), .B(\u_div/u_add_PartRem_2_16/n2 ), 
        .Y(\u_div/CryTmp[16][6] ) );
  XNOR2X1 U390 ( .A(\u_div/PartRem[17][3] ), .B(\u_div/PartRem[17][2] ), .Y(
        \u_div/SumTmp[16][3] ) );
  XNOR2X1 U391 ( .A(\u_div/PartRem[16][3] ), .B(\u_div/PartRem[16][2] ), .Y(
        \u_div/SumTmp[15][3] ) );
  OR2X1 U392 ( .A(\u_div/PartRem[15][5] ), .B(\u_div/u_add_PartRem_2_14/n2 ), 
        .Y(\u_div/CryTmp[14][6] ) );
  XNOR2X1 U393 ( .A(\u_div/PartRem[15][3] ), .B(\u_div/PartRem[15][2] ), .Y(
        \u_div/SumTmp[14][3] ) );
  OR2X1 U394 ( .A(\u_div/PartRem[14][5] ), .B(\u_div/u_add_PartRem_2_13/n2 ), 
        .Y(\u_div/CryTmp[13][6] ) );
  XNOR2X1 U395 ( .A(\u_div/PartRem[14][3] ), .B(\u_div/PartRem[14][2] ), .Y(
        \u_div/SumTmp[13][3] ) );
  OR2X1 U396 ( .A(\u_div/PartRem[13][5] ), .B(\u_div/u_add_PartRem_2_12/n2 ), 
        .Y(\u_div/CryTmp[12][6] ) );
  XNOR2X1 U397 ( .A(\u_div/PartRem[13][3] ), .B(\u_div/PartRem[13][2] ), .Y(
        \u_div/SumTmp[12][3] ) );
  OR2X1 U398 ( .A(\u_div/PartRem[13][2] ), .B(\u_div/PartRem[13][3] ), .Y(
        \u_div/u_add_PartRem_2_12/n3 ) );
  OR2X1 U399 ( .A(\u_div/PartRem[12][5] ), .B(\u_div/u_add_PartRem_2_11/n2 ), 
        .Y(\u_div/CryTmp[11][6] ) );
  XNOR2X1 U400 ( .A(\u_div/PartRem[12][3] ), .B(\u_div/PartRem[12][2] ), .Y(
        \u_div/SumTmp[11][3] ) );
  XNOR2X1 U401 ( .A(\u_div/PartRem[11][3] ), .B(\u_div/PartRem[11][2] ), .Y(
        \u_div/SumTmp[10][3] ) );
  XNOR2X1 U402 ( .A(\u_div/PartRem[10][3] ), .B(\u_div/PartRem[10][2] ), .Y(
        \u_div/SumTmp[9][3] ) );
  XNOR2X1 U403 ( .A(\u_div/PartRem[9][3] ), .B(\u_div/PartRem[9][2] ), .Y(
        \u_div/SumTmp[8][3] ) );
  XNOR2X1 U404 ( .A(\u_div/PartRem[8][3] ), .B(\u_div/PartRem[8][2] ), .Y(
        \u_div/SumTmp[7][3] ) );
  OR2X1 U405 ( .A(\u_div/PartRem[8][2] ), .B(\u_div/PartRem[8][3] ), .Y(
        \u_div/u_add_PartRem_2_7/n3 ) );
  XNOR2X1 U406 ( .A(\u_div/PartRem[7][3] ), .B(\u_div/PartRem[7][2] ), .Y(
        \u_div/SumTmp[6][3] ) );
  XNOR2X1 U407 ( .A(\u_div/PartRem[6][3] ), .B(\u_div/PartRem[6][2] ), .Y(
        \u_div/SumTmp[5][3] ) );
  XNOR2X1 U408 ( .A(\u_div/PartRem[5][3] ), .B(\u_div/PartRem[5][2] ), .Y(
        \u_div/SumTmp[4][3] ) );
  XNOR2X1 U409 ( .A(\u_div/PartRem[4][3] ), .B(\u_div/PartRem[4][2] ), .Y(
        \u_div/SumTmp[3][3] ) );
  XNOR2X1 U410 ( .A(\u_div/PartRem[3][3] ), .B(\u_div/PartRem[3][2] ), .Y(
        \u_div/SumTmp[2][3] ) );
  OR2X1 U411 ( .A(\u_div/PartRem[3][2] ), .B(\u_div/PartRem[3][3] ), .Y(
        \u_div/u_add_PartRem_2_2/n3 ) );
  OR2X1 U412 ( .A(\u_div/PartRem[2][5] ), .B(\u_div/u_add_PartRem_2_1/n2 ), 
        .Y(\u_div/CryTmp[1][6] ) );
  XNOR2X1 U413 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/PartRem[2][2] ), .Y(
        \u_div/SumTmp[1][3] ) );
  NAND2BX1 U414 ( .AN(\u_div/PartRem[1][3] ), .B(n1), .Y(n6) );
  XNOR2X1 U415 ( .A(\u_div/PartRem[63][0] ), .B(\u_div/PartRem[62][0] ), .Y(
        \u_div/SumTmp[59][3] ) );
  XOR2X1 U416 ( .A(\u_div/CryTmp[58][6] ), .B(n4), .Y(\u_div/QInv[58] ) );
  XOR2X1 U417 ( .A(\u_div/CryTmp[39][6] ), .B(n4), .Y(\u_div/QInv[39] ) );
  XOR2X1 U418 ( .A(\u_div/CryTmp[29][6] ), .B(n4), .Y(\u_div/QInv[29] ) );
  XOR2X1 U419 ( .A(\u_div/CryTmp[18][6] ), .B(n4), .Y(\u_div/QInv[18] ) );
  XOR2X1 U420 ( .A(\u_div/CryTmp[0][6] ), .B(n4), .Y(\u_div/QInv[0] ) );
endmodule


module GSIM_DW01_inc_7 ( A, SUM );
  input [63:0] A;
  output [63:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;

  NOR3BX1 U2 ( .AN(A[59]), .B(n1), .C(n24), .Y(n22) );
  NOR3BX1 U3 ( .AN(A[55]), .B(n2), .C(n30), .Y(n28) );
  NOR3BX1 U4 ( .AN(A[51]), .B(n3), .C(n34), .Y(n32) );
  NOR3BX1 U5 ( .AN(A[47]), .B(n4), .C(n38), .Y(n36) );
  NOR3BX1 U6 ( .AN(A[43]), .B(n5), .C(n42), .Y(n40) );
  NOR3BX1 U7 ( .AN(A[39]), .B(n6), .C(n46), .Y(n44) );
  NOR3BX1 U8 ( .AN(A[35]), .B(n7), .C(n52), .Y(n50) );
  NOR3BX1 U9 ( .AN(A[31]), .B(n8), .C(n56), .Y(n54) );
  NOR3BX1 U10 ( .AN(A[27]), .B(n9), .C(n60), .Y(n58) );
  NOR3BX1 U11 ( .AN(A[23]), .B(n10), .C(n64), .Y(n62) );
  NOR3BX1 U12 ( .AN(A[19]), .B(n11), .C(n68), .Y(n66) );
  NOR3BX1 U13 ( .AN(A[15]), .B(n12), .C(n72), .Y(n70) );
  NOR3BX1 U14 ( .AN(A[11]), .B(n13), .C(n76), .Y(n74) );
  NOR3BX1 U15 ( .AN(A[7]), .B(n14), .C(n19), .Y(n17) );
  NAND3X1 U16 ( .A(A[4]), .B(n26), .C(A[5]), .Y(n19) );
  NOR3BX1 U17 ( .AN(A[3]), .B(n15), .C(n48), .Y(n26) );
  NOR2XL U18 ( .A(n24), .B(n1), .Y(n27) );
  NAND2XL U19 ( .A(A[56]), .B(n28), .Y(n29) );
  NOR2XL U20 ( .A(n30), .B(n2), .Y(n31) );
  NAND2XL U21 ( .A(A[52]), .B(n32), .Y(n33) );
  NOR2XL U22 ( .A(n34), .B(n3), .Y(n35) );
  NAND2XL U23 ( .A(A[48]), .B(n36), .Y(n37) );
  NOR2XL U24 ( .A(n38), .B(n4), .Y(n39) );
  NAND2XL U25 ( .A(A[44]), .B(n40), .Y(n41) );
  NOR2XL U26 ( .A(n42), .B(n5), .Y(n43) );
  NAND2XL U27 ( .A(A[40]), .B(n44), .Y(n45) );
  NOR2XL U28 ( .A(n46), .B(n6), .Y(n49) );
  NAND2XL U29 ( .A(A[36]), .B(n50), .Y(n51) );
  NOR2XL U30 ( .A(n52), .B(n7), .Y(n53) );
  NAND2XL U31 ( .A(A[32]), .B(n54), .Y(n55) );
  NOR2XL U32 ( .A(n56), .B(n8), .Y(n57) );
  NAND2XL U33 ( .A(A[28]), .B(n58), .Y(n59) );
  NOR2XL U34 ( .A(n60), .B(n9), .Y(n61) );
  NAND2XL U35 ( .A(A[24]), .B(n62), .Y(n63) );
  NOR2XL U36 ( .A(n64), .B(n10), .Y(n65) );
  NAND2XL U37 ( .A(A[20]), .B(n66), .Y(n67) );
  NOR2XL U38 ( .A(n68), .B(n11), .Y(n69) );
  NAND2XL U39 ( .A(A[16]), .B(n70), .Y(n71) );
  NOR2XL U40 ( .A(n72), .B(n12), .Y(n73) );
  NAND2XL U41 ( .A(A[12]), .B(n74), .Y(n75) );
  NOR2XL U42 ( .A(n76), .B(n13), .Y(n77) );
  NAND2XL U43 ( .A(A[8]), .B(n17), .Y(n16) );
  NOR2XL U44 ( .A(n19), .B(n14), .Y(n18) );
  NAND2XL U45 ( .A(A[4]), .B(n26), .Y(n25) );
  XOR2XL U46 ( .A(A[60]), .B(n22), .Y(SUM[60]) );
  NAND2XL U47 ( .A(A[60]), .B(n22), .Y(n23) );
  NOR2XL U48 ( .A(n48), .B(n15), .Y(n47) );
  XOR2X1 U49 ( .A(A[63]), .B(n20), .Y(SUM[63]) );
  CLKINVX1 U50 ( .A(A[2]), .Y(n15) );
  CLKINVX1 U51 ( .A(A[42]), .Y(n5) );
  CLKINVX1 U52 ( .A(A[30]), .Y(n8) );
  CLKINVX1 U53 ( .A(A[26]), .Y(n9) );
  CLKINVX1 U54 ( .A(A[22]), .Y(n10) );
  CLKINVX1 U55 ( .A(A[18]), .Y(n11) );
  CLKINVX1 U56 ( .A(A[14]), .Y(n12) );
  CLKINVX1 U57 ( .A(A[10]), .Y(n13) );
  CLKINVX1 U58 ( .A(A[6]), .Y(n14) );
  CLKINVX1 U59 ( .A(A[58]), .Y(n1) );
  CLKINVX1 U60 ( .A(A[38]), .Y(n6) );
  CLKINVX1 U61 ( .A(A[34]), .Y(n7) );
  CLKINVX1 U62 ( .A(A[54]), .Y(n2) );
  CLKINVX1 U63 ( .A(A[50]), .Y(n3) );
  CLKINVX1 U64 ( .A(A[46]), .Y(n4) );
  XNOR2X1 U65 ( .A(A[9]), .B(n16), .Y(SUM[9]) );
  XOR2X1 U66 ( .A(A[8]), .B(n17), .Y(SUM[8]) );
  XOR2X1 U67 ( .A(A[7]), .B(n18), .Y(SUM[7]) );
  XOR2X1 U68 ( .A(n14), .B(n19), .Y(SUM[6]) );
  NOR2BX1 U69 ( .AN(A[62]), .B(n21), .Y(n20) );
  XNOR2X1 U70 ( .A(A[62]), .B(n21), .Y(SUM[62]) );
  NAND3X1 U71 ( .A(A[60]), .B(n22), .C(A[61]), .Y(n21) );
  XNOR2X1 U72 ( .A(A[61]), .B(n23), .Y(SUM[61]) );
  XNOR2X1 U73 ( .A(A[5]), .B(n25), .Y(SUM[5]) );
  XOR2X1 U74 ( .A(A[59]), .B(n27), .Y(SUM[59]) );
  XOR2X1 U75 ( .A(n1), .B(n24), .Y(SUM[58]) );
  NAND3X1 U76 ( .A(A[56]), .B(n28), .C(A[57]), .Y(n24) );
  XNOR2X1 U77 ( .A(A[57]), .B(n29), .Y(SUM[57]) );
  XOR2X1 U78 ( .A(A[56]), .B(n28), .Y(SUM[56]) );
  XOR2X1 U79 ( .A(A[55]), .B(n31), .Y(SUM[55]) );
  XOR2X1 U80 ( .A(n2), .B(n30), .Y(SUM[54]) );
  NAND3X1 U81 ( .A(A[52]), .B(n32), .C(A[53]), .Y(n30) );
  XNOR2X1 U82 ( .A(A[53]), .B(n33), .Y(SUM[53]) );
  XOR2X1 U83 ( .A(A[52]), .B(n32), .Y(SUM[52]) );
  XOR2X1 U84 ( .A(A[51]), .B(n35), .Y(SUM[51]) );
  XOR2X1 U85 ( .A(n3), .B(n34), .Y(SUM[50]) );
  NAND3X1 U86 ( .A(A[48]), .B(n36), .C(A[49]), .Y(n34) );
  XOR2X1 U87 ( .A(A[4]), .B(n26), .Y(SUM[4]) );
  XNOR2X1 U88 ( .A(A[49]), .B(n37), .Y(SUM[49]) );
  XOR2X1 U89 ( .A(A[48]), .B(n36), .Y(SUM[48]) );
  XOR2X1 U90 ( .A(A[47]), .B(n39), .Y(SUM[47]) );
  XOR2X1 U91 ( .A(n4), .B(n38), .Y(SUM[46]) );
  NAND3X1 U92 ( .A(A[44]), .B(n40), .C(A[45]), .Y(n38) );
  XNOR2X1 U93 ( .A(A[45]), .B(n41), .Y(SUM[45]) );
  XOR2X1 U94 ( .A(A[44]), .B(n40), .Y(SUM[44]) );
  XOR2X1 U95 ( .A(A[43]), .B(n43), .Y(SUM[43]) );
  XOR2X1 U96 ( .A(n5), .B(n42), .Y(SUM[42]) );
  NAND3X1 U97 ( .A(A[40]), .B(n44), .C(A[41]), .Y(n42) );
  XNOR2X1 U98 ( .A(A[41]), .B(n45), .Y(SUM[41]) );
  XOR2X1 U99 ( .A(A[40]), .B(n44), .Y(SUM[40]) );
  XOR2X1 U100 ( .A(A[3]), .B(n47), .Y(SUM[3]) );
  XOR2X1 U101 ( .A(A[39]), .B(n49), .Y(SUM[39]) );
  XOR2X1 U102 ( .A(n6), .B(n46), .Y(SUM[38]) );
  NAND3X1 U103 ( .A(A[36]), .B(n50), .C(A[37]), .Y(n46) );
  XNOR2X1 U104 ( .A(A[37]), .B(n51), .Y(SUM[37]) );
  XOR2X1 U105 ( .A(A[36]), .B(n50), .Y(SUM[36]) );
  XOR2X1 U106 ( .A(A[35]), .B(n53), .Y(SUM[35]) );
  XOR2X1 U107 ( .A(n7), .B(n52), .Y(SUM[34]) );
  NAND3X1 U108 ( .A(A[32]), .B(n54), .C(A[33]), .Y(n52) );
  XNOR2X1 U109 ( .A(A[33]), .B(n55), .Y(SUM[33]) );
  XOR2X1 U110 ( .A(A[32]), .B(n54), .Y(SUM[32]) );
  XOR2X1 U111 ( .A(A[31]), .B(n57), .Y(SUM[31]) );
  XOR2X1 U112 ( .A(n8), .B(n56), .Y(SUM[30]) );
  NAND3X1 U113 ( .A(A[28]), .B(n58), .C(A[29]), .Y(n56) );
  XOR2X1 U114 ( .A(n15), .B(n48), .Y(SUM[2]) );
  XNOR2X1 U115 ( .A(A[29]), .B(n59), .Y(SUM[29]) );
  XOR2X1 U116 ( .A(A[28]), .B(n58), .Y(SUM[28]) );
  XOR2X1 U117 ( .A(A[27]), .B(n61), .Y(SUM[27]) );
  XOR2X1 U118 ( .A(n9), .B(n60), .Y(SUM[26]) );
  NAND3X1 U119 ( .A(A[24]), .B(n62), .C(A[25]), .Y(n60) );
  XNOR2X1 U120 ( .A(A[25]), .B(n63), .Y(SUM[25]) );
  XOR2X1 U121 ( .A(A[24]), .B(n62), .Y(SUM[24]) );
  XOR2X1 U122 ( .A(A[23]), .B(n65), .Y(SUM[23]) );
  XOR2X1 U123 ( .A(n10), .B(n64), .Y(SUM[22]) );
  NAND3X1 U124 ( .A(A[20]), .B(n66), .C(A[21]), .Y(n64) );
  XNOR2X1 U125 ( .A(A[21]), .B(n67), .Y(SUM[21]) );
  XOR2X1 U126 ( .A(A[20]), .B(n66), .Y(SUM[20]) );
  XOR2X1 U127 ( .A(A[19]), .B(n69), .Y(SUM[19]) );
  XOR2X1 U128 ( .A(n11), .B(n68), .Y(SUM[18]) );
  NAND3X1 U129 ( .A(A[16]), .B(n70), .C(A[17]), .Y(n68) );
  XNOR2X1 U130 ( .A(A[17]), .B(n71), .Y(SUM[17]) );
  XOR2X1 U131 ( .A(A[16]), .B(n70), .Y(SUM[16]) );
  XOR2X1 U132 ( .A(A[15]), .B(n73), .Y(SUM[15]) );
  XOR2X1 U133 ( .A(n12), .B(n72), .Y(SUM[14]) );
  NAND3X1 U134 ( .A(A[12]), .B(n74), .C(A[13]), .Y(n72) );
  XNOR2X1 U135 ( .A(A[13]), .B(n75), .Y(SUM[13]) );
  XOR2X1 U136 ( .A(A[12]), .B(n74), .Y(SUM[12]) );
  XOR2X1 U137 ( .A(A[11]), .B(n77), .Y(SUM[11]) );
  XOR2X1 U138 ( .A(n13), .B(n76), .Y(SUM[10]) );
  NAND3X1 U139 ( .A(A[8]), .B(n17), .C(A[9]), .Y(n76) );
  NAND2X1 U140 ( .A(A[1]), .B(A[0]), .Y(n48) );
endmodule


module GSIM_DW01_absval_5 ( A, ABSVAL );
  input [63:0] A;
  output [63:0] ABSVAL;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68;
  wire   [63:0] AMUX1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  GSIM_DW01_inc_7 NEG ( .A({n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
        n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
        n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
        n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
        n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68}), .SUM({
        AMUX1[63:2], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1}) );
  CLKINVX1 U1 ( .A(A[61]), .Y(n7) );
  CLKMX2X3 U2 ( .A(A[61]), .B(AMUX1[61]), .S0(n4), .Y(ABSVAL[61]) );
  CLKINVX1 U3 ( .A(A[3]), .Y(n65) );
  INVX3 U4 ( .A(n5), .Y(n4) );
  INVX3 U5 ( .A(n5), .Y(n3) );
  INVX3 U6 ( .A(n5), .Y(n2) );
  INVX3 U7 ( .A(n5), .Y(n1) );
  CLKINVX1 U8 ( .A(A[63]), .Y(n5) );
  AND2X2 U9 ( .A(AMUX1[63]), .B(n4), .Y(ABSVAL[63]) );
  CLKINVX1 U10 ( .A(A[2]), .Y(n66) );
  CLKINVX1 U11 ( .A(A[4]), .Y(n64) );
  CLKINVX1 U12 ( .A(A[42]), .Y(n26) );
  CLKINVX1 U13 ( .A(A[30]), .Y(n38) );
  CLKINVX1 U14 ( .A(A[26]), .Y(n42) );
  CLKINVX1 U15 ( .A(A[22]), .Y(n46) );
  CLKINVX1 U16 ( .A(A[18]), .Y(n50) );
  CLKINVX1 U17 ( .A(A[14]), .Y(n54) );
  CLKINVX1 U18 ( .A(A[10]), .Y(n58) );
  CLKINVX1 U19 ( .A(A[6]), .Y(n62) );
  CLKINVX1 U20 ( .A(A[29]), .Y(n39) );
  CLKINVX1 U21 ( .A(A[21]), .Y(n47) );
  CLKINVX1 U22 ( .A(A[17]), .Y(n51) );
  CLKINVX1 U23 ( .A(A[13]), .Y(n55) );
  CLKINVX1 U24 ( .A(A[9]), .Y(n59) );
  CLKINVX1 U25 ( .A(A[5]), .Y(n63) );
  CLKINVX1 U26 ( .A(A[51]), .Y(n17) );
  CLKINVX1 U27 ( .A(A[47]), .Y(n21) );
  CLKINVX1 U28 ( .A(A[43]), .Y(n25) );
  CLKINVX1 U29 ( .A(A[39]), .Y(n29) );
  CLKINVX1 U30 ( .A(A[35]), .Y(n33) );
  CLKINVX1 U31 ( .A(A[31]), .Y(n37) );
  CLKINVX1 U32 ( .A(A[27]), .Y(n41) );
  CLKINVX1 U33 ( .A(A[23]), .Y(n45) );
  CLKINVX1 U34 ( .A(A[19]), .Y(n49) );
  CLKINVX1 U35 ( .A(A[15]), .Y(n53) );
  CLKINVX1 U36 ( .A(A[11]), .Y(n57) );
  CLKINVX1 U37 ( .A(A[7]), .Y(n61) );
  CLKINVX1 U38 ( .A(A[52]), .Y(n16) );
  CLKINVX1 U39 ( .A(A[48]), .Y(n20) );
  CLKINVX1 U40 ( .A(A[40]), .Y(n28) );
  CLKINVX1 U41 ( .A(A[36]), .Y(n32) );
  CLKINVX1 U42 ( .A(A[32]), .Y(n36) );
  CLKINVX1 U43 ( .A(A[28]), .Y(n40) );
  CLKINVX1 U44 ( .A(A[24]), .Y(n44) );
  CLKINVX1 U45 ( .A(A[20]), .Y(n48) );
  CLKINVX1 U46 ( .A(A[16]), .Y(n52) );
  CLKINVX1 U47 ( .A(A[12]), .Y(n56) );
  CLKINVX1 U48 ( .A(A[8]), .Y(n60) );
  CLKINVX1 U49 ( .A(A[58]), .Y(n10) );
  CLKINVX1 U50 ( .A(A[38]), .Y(n30) );
  CLKINVX1 U51 ( .A(A[34]), .Y(n34) );
  CLKINVX1 U52 ( .A(A[57]), .Y(n11) );
  CLKINVX1 U53 ( .A(A[53]), .Y(n15) );
  CLKINVX1 U54 ( .A(A[49]), .Y(n19) );
  CLKINVX1 U55 ( .A(A[45]), .Y(n23) );
  CLKINVX1 U56 ( .A(A[41]), .Y(n27) );
  CLKINVX1 U57 ( .A(A[37]), .Y(n31) );
  CLKINVX1 U58 ( .A(A[33]), .Y(n35) );
  CLKINVX1 U59 ( .A(A[25]), .Y(n43) );
  CLKINVX1 U60 ( .A(A[62]), .Y(n6) );
  CLKINVX1 U61 ( .A(A[59]), .Y(n9) );
  CLKINVX1 U62 ( .A(A[55]), .Y(n13) );
  CLKINVX1 U63 ( .A(A[54]), .Y(n14) );
  CLKINVX1 U64 ( .A(A[50]), .Y(n18) );
  CLKINVX1 U65 ( .A(A[46]), .Y(n22) );
  CLKINVX1 U66 ( .A(A[60]), .Y(n8) );
  CLKINVX1 U67 ( .A(A[56]), .Y(n12) );
  CLKINVX1 U68 ( .A(A[44]), .Y(n24) );
  CLKINVX1 U69 ( .A(A[0]), .Y(n68) );
  CLKINVX1 U70 ( .A(A[1]), .Y(n67) );
  CLKMX2X2 U71 ( .A(A[9]), .B(AMUX1[9]), .S0(n3), .Y(ABSVAL[9]) );
  CLKMX2X2 U72 ( .A(A[8]), .B(AMUX1[8]), .S0(n4), .Y(ABSVAL[8]) );
  CLKMX2X2 U73 ( .A(A[7]), .B(AMUX1[7]), .S0(n4), .Y(ABSVAL[7]) );
  CLKMX2X2 U74 ( .A(A[6]), .B(AMUX1[6]), .S0(n4), .Y(ABSVAL[6]) );
  CLKMX2X2 U75 ( .A(A[62]), .B(AMUX1[62]), .S0(n4), .Y(ABSVAL[62]) );
  CLKMX2X2 U76 ( .A(A[60]), .B(AMUX1[60]), .S0(n4), .Y(ABSVAL[60]) );
  CLKMX2X2 U77 ( .A(A[5]), .B(AMUX1[5]), .S0(n4), .Y(ABSVAL[5]) );
  CLKMX2X2 U78 ( .A(A[59]), .B(AMUX1[59]), .S0(n4), .Y(ABSVAL[59]) );
  CLKMX2X2 U79 ( .A(A[58]), .B(AMUX1[58]), .S0(n4), .Y(ABSVAL[58]) );
  CLKMX2X2 U80 ( .A(A[57]), .B(AMUX1[57]), .S0(n4), .Y(ABSVAL[57]) );
  CLKMX2X2 U81 ( .A(A[56]), .B(AMUX1[56]), .S0(n3), .Y(ABSVAL[56]) );
  CLKMX2X2 U82 ( .A(A[55]), .B(AMUX1[55]), .S0(n3), .Y(ABSVAL[55]) );
  CLKMX2X2 U83 ( .A(A[54]), .B(AMUX1[54]), .S0(n3), .Y(ABSVAL[54]) );
  CLKMX2X2 U84 ( .A(A[53]), .B(AMUX1[53]), .S0(n3), .Y(ABSVAL[53]) );
  CLKMX2X2 U85 ( .A(A[52]), .B(AMUX1[52]), .S0(n3), .Y(ABSVAL[52]) );
  CLKMX2X2 U86 ( .A(A[51]), .B(AMUX1[51]), .S0(n3), .Y(ABSVAL[51]) );
  CLKMX2X2 U87 ( .A(A[50]), .B(AMUX1[50]), .S0(n3), .Y(ABSVAL[50]) );
  CLKMX2X2 U88 ( .A(A[4]), .B(AMUX1[4]), .S0(n3), .Y(ABSVAL[4]) );
  CLKMX2X2 U89 ( .A(A[49]), .B(AMUX1[49]), .S0(n3), .Y(ABSVAL[49]) );
  CLKMX2X2 U90 ( .A(A[48]), .B(AMUX1[48]), .S0(n3), .Y(ABSVAL[48]) );
  CLKMX2X2 U91 ( .A(A[47]), .B(AMUX1[47]), .S0(n3), .Y(ABSVAL[47]) );
  CLKMX2X2 U92 ( .A(A[46]), .B(AMUX1[46]), .S0(n3), .Y(ABSVAL[46]) );
  CLKMX2X2 U93 ( .A(A[45]), .B(AMUX1[45]), .S0(n3), .Y(ABSVAL[45]) );
  CLKMX2X2 U94 ( .A(A[44]), .B(AMUX1[44]), .S0(n2), .Y(ABSVAL[44]) );
  CLKMX2X2 U95 ( .A(A[43]), .B(AMUX1[43]), .S0(n2), .Y(ABSVAL[43]) );
  CLKMX2X2 U96 ( .A(A[42]), .B(AMUX1[42]), .S0(n2), .Y(ABSVAL[42]) );
  CLKMX2X2 U97 ( .A(A[41]), .B(AMUX1[41]), .S0(n2), .Y(ABSVAL[41]) );
  CLKMX2X2 U98 ( .A(A[40]), .B(AMUX1[40]), .S0(n2), .Y(ABSVAL[40]) );
  CLKMX2X2 U99 ( .A(A[3]), .B(AMUX1[3]), .S0(n2), .Y(ABSVAL[3]) );
  CLKMX2X2 U100 ( .A(A[39]), .B(AMUX1[39]), .S0(n2), .Y(ABSVAL[39]) );
  CLKMX2X2 U101 ( .A(A[38]), .B(AMUX1[38]), .S0(n2), .Y(ABSVAL[38]) );
  CLKMX2X2 U102 ( .A(A[37]), .B(AMUX1[37]), .S0(n2), .Y(ABSVAL[37]) );
  CLKMX2X2 U103 ( .A(A[36]), .B(AMUX1[36]), .S0(n2), .Y(ABSVAL[36]) );
  CLKMX2X2 U104 ( .A(A[35]), .B(AMUX1[35]), .S0(n2), .Y(ABSVAL[35]) );
  CLKMX2X2 U105 ( .A(A[34]), .B(AMUX1[34]), .S0(n2), .Y(ABSVAL[34]) );
  CLKMX2X2 U106 ( .A(A[33]), .B(AMUX1[33]), .S0(n1), .Y(ABSVAL[33]) );
  CLKMX2X2 U107 ( .A(A[32]), .B(AMUX1[32]), .S0(n1), .Y(ABSVAL[32]) );
  CLKMX2X2 U108 ( .A(A[31]), .B(AMUX1[31]), .S0(n1), .Y(ABSVAL[31]) );
  CLKMX2X2 U109 ( .A(A[30]), .B(AMUX1[30]), .S0(n1), .Y(ABSVAL[30]) );
  CLKMX2X2 U110 ( .A(A[2]), .B(AMUX1[2]), .S0(n1), .Y(ABSVAL[2]) );
  CLKMX2X2 U111 ( .A(A[29]), .B(AMUX1[29]), .S0(n1), .Y(ABSVAL[29]) );
  CLKMX2X2 U112 ( .A(A[28]), .B(AMUX1[28]), .S0(n1), .Y(ABSVAL[28]) );
  CLKMX2X2 U113 ( .A(A[27]), .B(AMUX1[27]), .S0(n1), .Y(ABSVAL[27]) );
  CLKMX2X2 U114 ( .A(A[26]), .B(AMUX1[26]), .S0(n1), .Y(ABSVAL[26]) );
  CLKMX2X2 U115 ( .A(A[25]), .B(AMUX1[25]), .S0(n1), .Y(ABSVAL[25]) );
  CLKMX2X2 U116 ( .A(A[24]), .B(AMUX1[24]), .S0(n1), .Y(ABSVAL[24]) );
  CLKMX2X2 U117 ( .A(A[23]), .B(AMUX1[23]), .S0(n1), .Y(ABSVAL[23]) );
  CLKMX2X2 U118 ( .A(A[22]), .B(AMUX1[22]), .S0(n1), .Y(ABSVAL[22]) );
  CLKMX2X2 U119 ( .A(A[21]), .B(AMUX1[21]), .S0(n1), .Y(ABSVAL[21]) );
  CLKMX2X2 U120 ( .A(A[20]), .B(AMUX1[20]), .S0(n1), .Y(ABSVAL[20]) );
  CLKMX2X2 U121 ( .A(A[19]), .B(AMUX1[19]), .S0(n1), .Y(ABSVAL[19]) );
  CLKMX2X2 U122 ( .A(A[18]), .B(AMUX1[18]), .S0(n1), .Y(ABSVAL[18]) );
  CLKMX2X2 U123 ( .A(A[17]), .B(AMUX1[17]), .S0(n2), .Y(ABSVAL[17]) );
  CLKMX2X2 U124 ( .A(A[16]), .B(AMUX1[16]), .S0(n2), .Y(ABSVAL[16]) );
  CLKMX2X2 U125 ( .A(A[15]), .B(AMUX1[15]), .S0(n2), .Y(ABSVAL[15]) );
  CLKMX2X2 U126 ( .A(A[14]), .B(AMUX1[14]), .S0(n2), .Y(ABSVAL[14]) );
  CLKMX2X2 U127 ( .A(A[13]), .B(AMUX1[13]), .S0(n3), .Y(ABSVAL[13]) );
  CLKMX2X2 U128 ( .A(A[12]), .B(AMUX1[12]), .S0(n3), .Y(ABSVAL[12]) );
  CLKMX2X2 U129 ( .A(A[11]), .B(AMUX1[11]), .S0(n3), .Y(ABSVAL[11]) );
  CLKMX2X2 U130 ( .A(A[10]), .B(AMUX1[10]), .S0(n2), .Y(ABSVAL[10]) );
endmodule


module GSIM_DW_inc_5 ( carry_in, a, carry_out, sum );
  input [63:0] a;
  output [63:0] sum;
  input carry_in;
  output carry_out;
  wire   \sum[63] , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63;
  assign sum[62] = \sum[63] ;
  assign sum[61] = \sum[63] ;
  assign sum[63] = \sum[63] ;

  ADDHXL U20 ( .A(a[46]), .B(n18), .CO(n17), .S(sum[46]) );
  ADDHXL U38 ( .A(a[28]), .B(n36), .CO(n35), .S(sum[28]) );
  ADDHXL U41 ( .A(a[25]), .B(n39), .CO(n38), .S(sum[25]) );
  ADDHXL U60 ( .A(a[6]), .B(n58), .CO(n57), .S(sum[6]) );
  ADDHX2 U70 ( .A(a[29]), .B(n35), .CO(n34), .S(sum[29]) );
  ADDHX2 U71 ( .A(a[41]), .B(n23), .CO(n22), .S(sum[41]) );
  ADDHX2 U72 ( .A(a[31]), .B(n33), .CO(n32), .S(sum[31]) );
  ADDHX2 U73 ( .A(a[12]), .B(n52), .CO(n51), .S(sum[12]) );
  ADDHX2 U74 ( .A(a[14]), .B(n50), .CO(n49), .S(sum[14]) );
  ADDHX2 U75 ( .A(a[39]), .B(n25), .CO(n24), .S(sum[39]) );
  ADDHX2 U76 ( .A(a[35]), .B(n29), .CO(n28), .S(sum[35]) );
  ADDHX1 U77 ( .A(a[7]), .B(n57), .CO(n56), .S(sum[7]) );
  ADDHX2 U78 ( .A(a[16]), .B(n48), .CO(n47), .S(sum[16]) );
  ADDHX1 U79 ( .A(carry_in), .B(a[0]), .CO(n63), .S(sum[0]) );
  ADDHXL U80 ( .A(a[36]), .B(n28), .CO(n27), .S(sum[36]) );
  ADDHXL U81 ( .A(a[17]), .B(n47), .CO(n46), .S(sum[17]) );
  ADDHXL U82 ( .A(a[8]), .B(n56), .CO(n55), .S(sum[8]) );
  ADDHX2 U83 ( .A(a[52]), .B(n12), .CO(n11), .S(sum[52]) );
  ADDHX2 U84 ( .A(a[40]), .B(n24), .CO(n23), .S(sum[40]) );
  ADDHX2 U85 ( .A(a[13]), .B(n51), .CO(n50), .S(sum[13]) );
  ADDHX2 U86 ( .A(a[30]), .B(n34), .CO(n33), .S(sum[30]) );
  ADDHX2 U87 ( .A(a[15]), .B(n49), .CO(n48), .S(sum[15]) );
  ADDHX2 U88 ( .A(a[56]), .B(n8), .CO(n7), .S(sum[56]) );
  ADDHX2 U89 ( .A(a[9]), .B(n55), .CO(n54), .S(sum[9]) );
  ADDHX2 U90 ( .A(a[42]), .B(n22), .CO(n21), .S(sum[42]) );
  ADDHX2 U91 ( .A(a[37]), .B(n27), .CO(n26), .S(sum[37]) );
  ADDHX2 U92 ( .A(a[32]), .B(n32), .CO(n31), .S(sum[32]) );
  XOR2X4 U93 ( .A(n4), .B(a[60]), .Y(sum[60]) );
  NOR2BX1 U94 ( .AN(a[60]), .B(n4), .Y(\sum[63] ) );
  ADDHX2 U95 ( .A(a[58]), .B(n6), .CO(n5), .S(sum[58]) );
  ADDHX1 U96 ( .A(a[55]), .B(n9), .CO(n8), .S(sum[55]) );
  ADDHX1 U97 ( .A(a[47]), .B(n17), .CO(n16), .S(sum[47]) );
  ADDHX1 U98 ( .A(a[44]), .B(n20), .CO(n19), .S(sum[44]) );
  ADDHX1 U99 ( .A(a[34]), .B(n30), .CO(n29), .S(sum[34]) );
  ADDHX1 U100 ( .A(a[11]), .B(n53), .CO(n52), .S(sum[11]) );
  ADDHX1 U101 ( .A(a[26]), .B(n38), .CO(n37), .S(sum[26]) );
  ADDHX1 U102 ( .A(a[23]), .B(n41), .CO(n40), .S(sum[23]) );
  ADDHX1 U103 ( .A(a[18]), .B(n46), .CO(n45), .S(sum[18]) );
  ADDHX1 U104 ( .A(a[5]), .B(n59), .CO(n58), .S(sum[5]) );
  ADDHX1 U105 ( .A(a[4]), .B(n60), .CO(n59), .S(sum[4]) );
  ADDHX1 U106 ( .A(a[1]), .B(n63), .CO(n62), .S(sum[1]) );
  ADDHX1 U107 ( .A(a[53]), .B(n11), .CO(n10), .S(sum[53]) );
  ADDHX1 U108 ( .A(a[50]), .B(n14), .CO(n13), .S(sum[50]) );
  ADDHX1 U109 ( .A(a[45]), .B(n19), .CO(n18), .S(sum[45]) );
  ADDHX1 U110 ( .A(a[48]), .B(n16), .CO(n15), .S(sum[48]) );
  ADDHX1 U111 ( .A(a[27]), .B(n37), .CO(n36), .S(sum[27]) );
  ADDHX1 U112 ( .A(a[24]), .B(n40), .CO(n39), .S(sum[24]) );
  ADDHX1 U113 ( .A(a[21]), .B(n43), .CO(n42), .S(sum[21]) );
  ADDHX1 U114 ( .A(a[19]), .B(n45), .CO(n44), .S(sum[19]) );
  ADDHX1 U115 ( .A(a[3]), .B(n61), .CO(n60), .S(sum[3]) );
  ADDHX1 U116 ( .A(a[2]), .B(n62), .CO(n61), .S(sum[2]) );
  ADDHXL U117 ( .A(a[59]), .B(n5), .CO(n4), .S(sum[59]) );
  ADDHXL U118 ( .A(a[10]), .B(n54), .CO(n53), .S(sum[10]) );
  ADDHXL U119 ( .A(a[20]), .B(n44), .CO(n43), .S(sum[20]) );
  ADDHXL U120 ( .A(a[22]), .B(n42), .CO(n41), .S(sum[22]) );
  ADDHXL U121 ( .A(a[57]), .B(n7), .CO(n6), .S(sum[57]) );
  ADDHXL U122 ( .A(a[51]), .B(n13), .CO(n12), .S(sum[51]) );
  ADDHXL U123 ( .A(a[49]), .B(n15), .CO(n14), .S(sum[49]) );
  ADDHXL U124 ( .A(a[54]), .B(n10), .CO(n9), .S(sum[54]) );
  ADDHXL U125 ( .A(a[33]), .B(n31), .CO(n30), .S(sum[33]) );
  ADDHXL U126 ( .A(a[43]), .B(n21), .CO(n20), .S(sum[43]) );
  ADDHXL U127 ( .A(a[38]), .B(n26), .CO(n25), .S(sum[38]) );
endmodule


module GSIM_DW_div_tc_5 ( a, b, quotient, remainder, divide_by_0 );
  input [63:0] a;
  input [5:0] b;
  output [63:0] quotient;
  output [5:0] remainder;
  output divide_by_0;
  wire   \u_div/QInv[63] , \u_div/QInv[59] , \u_div/QInv[58] ,
         \u_div/QInv[57] , \u_div/QInv[56] , \u_div/QInv[55] ,
         \u_div/QInv[54] , \u_div/QInv[53] , \u_div/QInv[52] ,
         \u_div/QInv[51] , \u_div/QInv[50] , \u_div/QInv[49] ,
         \u_div/QInv[48] , \u_div/QInv[47] , \u_div/QInv[46] ,
         \u_div/QInv[45] , \u_div/QInv[44] , \u_div/QInv[43] ,
         \u_div/QInv[42] , \u_div/QInv[41] , \u_div/QInv[40] ,
         \u_div/QInv[39] , \u_div/QInv[38] , \u_div/QInv[37] ,
         \u_div/QInv[36] , \u_div/QInv[35] , \u_div/QInv[34] ,
         \u_div/QInv[33] , \u_div/QInv[32] , \u_div/QInv[31] ,
         \u_div/QInv[30] , \u_div/QInv[29] , \u_div/QInv[28] ,
         \u_div/QInv[27] , \u_div/QInv[26] , \u_div/QInv[25] ,
         \u_div/QInv[24] , \u_div/QInv[23] , \u_div/QInv[22] ,
         \u_div/QInv[21] , \u_div/QInv[20] , \u_div/QInv[19] ,
         \u_div/QInv[18] , \u_div/QInv[17] , \u_div/QInv[16] ,
         \u_div/QInv[15] , \u_div/QInv[14] , \u_div/QInv[13] ,
         \u_div/QInv[12] , \u_div/QInv[11] , \u_div/QInv[10] , \u_div/QInv[9] ,
         \u_div/QInv[8] , \u_div/QInv[7] , \u_div/QInv[6] , \u_div/QInv[5] ,
         \u_div/QInv[4] , \u_div/QInv[3] , \u_div/QInv[2] , \u_div/QInv[1] ,
         \u_div/QInv[0] , \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] ,
         \u_div/SumTmp[1][3] , \u_div/SumTmp[1][4] , \u_div/SumTmp[2][1] ,
         \u_div/SumTmp[2][2] , \u_div/SumTmp[2][3] , \u_div/SumTmp[2][4] ,
         \u_div/SumTmp[3][1] , \u_div/SumTmp[3][2] , \u_div/SumTmp[3][3] ,
         \u_div/SumTmp[3][4] , \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] ,
         \u_div/SumTmp[4][3] , \u_div/SumTmp[4][4] , \u_div/SumTmp[5][1] ,
         \u_div/SumTmp[5][2] , \u_div/SumTmp[5][3] , \u_div/SumTmp[5][4] ,
         \u_div/SumTmp[6][1] , \u_div/SumTmp[6][2] , \u_div/SumTmp[6][3] ,
         \u_div/SumTmp[6][4] , \u_div/SumTmp[7][1] , \u_div/SumTmp[7][2] ,
         \u_div/SumTmp[7][3] , \u_div/SumTmp[7][4] , \u_div/SumTmp[8][1] ,
         \u_div/SumTmp[8][2] , \u_div/SumTmp[8][3] , \u_div/SumTmp[8][4] ,
         \u_div/SumTmp[9][1] , \u_div/SumTmp[9][2] , \u_div/SumTmp[9][3] ,
         \u_div/SumTmp[9][4] , \u_div/SumTmp[10][1] , \u_div/SumTmp[10][2] ,
         \u_div/SumTmp[10][3] , \u_div/SumTmp[10][4] , \u_div/SumTmp[11][1] ,
         \u_div/SumTmp[11][2] , \u_div/SumTmp[11][3] , \u_div/SumTmp[11][4] ,
         \u_div/SumTmp[12][1] , \u_div/SumTmp[12][2] , \u_div/SumTmp[12][3] ,
         \u_div/SumTmp[12][4] , \u_div/SumTmp[13][1] , \u_div/SumTmp[13][2] ,
         \u_div/SumTmp[13][3] , \u_div/SumTmp[13][4] , \u_div/SumTmp[14][1] ,
         \u_div/SumTmp[14][2] , \u_div/SumTmp[14][3] , \u_div/SumTmp[14][4] ,
         \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] , \u_div/SumTmp[15][3] ,
         \u_div/SumTmp[15][4] , \u_div/SumTmp[16][1] , \u_div/SumTmp[16][2] ,
         \u_div/SumTmp[16][3] , \u_div/SumTmp[16][4] , \u_div/SumTmp[17][1] ,
         \u_div/SumTmp[17][2] , \u_div/SumTmp[17][3] , \u_div/SumTmp[17][4] ,
         \u_div/SumTmp[18][1] , \u_div/SumTmp[18][2] , \u_div/SumTmp[18][3] ,
         \u_div/SumTmp[18][4] , \u_div/SumTmp[19][1] , \u_div/SumTmp[19][2] ,
         \u_div/SumTmp[19][3] , \u_div/SumTmp[19][4] , \u_div/SumTmp[20][1] ,
         \u_div/SumTmp[20][2] , \u_div/SumTmp[20][3] , \u_div/SumTmp[20][4] ,
         \u_div/SumTmp[21][1] , \u_div/SumTmp[21][2] , \u_div/SumTmp[21][3] ,
         \u_div/SumTmp[21][4] , \u_div/SumTmp[22][1] , \u_div/SumTmp[22][2] ,
         \u_div/SumTmp[22][3] , \u_div/SumTmp[22][4] , \u_div/SumTmp[23][1] ,
         \u_div/SumTmp[23][2] , \u_div/SumTmp[23][3] , \u_div/SumTmp[23][4] ,
         \u_div/SumTmp[24][1] , \u_div/SumTmp[24][2] , \u_div/SumTmp[24][3] ,
         \u_div/SumTmp[24][4] , \u_div/SumTmp[25][1] , \u_div/SumTmp[25][2] ,
         \u_div/SumTmp[25][3] , \u_div/SumTmp[25][4] , \u_div/SumTmp[26][1] ,
         \u_div/SumTmp[26][2] , \u_div/SumTmp[26][3] , \u_div/SumTmp[26][4] ,
         \u_div/SumTmp[27][1] , \u_div/SumTmp[27][2] , \u_div/SumTmp[27][3] ,
         \u_div/SumTmp[27][4] , \u_div/SumTmp[28][1] , \u_div/SumTmp[28][2] ,
         \u_div/SumTmp[28][3] , \u_div/SumTmp[28][4] , \u_div/SumTmp[29][1] ,
         \u_div/SumTmp[29][2] , \u_div/SumTmp[29][3] , \u_div/SumTmp[29][4] ,
         \u_div/SumTmp[30][1] , \u_div/SumTmp[30][2] , \u_div/SumTmp[30][3] ,
         \u_div/SumTmp[30][4] , \u_div/SumTmp[31][1] , \u_div/SumTmp[31][2] ,
         \u_div/SumTmp[31][3] , \u_div/SumTmp[31][4] , \u_div/SumTmp[32][1] ,
         \u_div/SumTmp[32][2] , \u_div/SumTmp[32][3] , \u_div/SumTmp[32][4] ,
         \u_div/SumTmp[33][1] , \u_div/SumTmp[33][2] , \u_div/SumTmp[33][3] ,
         \u_div/SumTmp[33][4] , \u_div/SumTmp[34][1] , \u_div/SumTmp[34][2] ,
         \u_div/SumTmp[34][3] , \u_div/SumTmp[34][4] , \u_div/SumTmp[35][1] ,
         \u_div/SumTmp[35][2] , \u_div/SumTmp[35][3] , \u_div/SumTmp[35][4] ,
         \u_div/SumTmp[36][1] , \u_div/SumTmp[36][2] , \u_div/SumTmp[36][3] ,
         \u_div/SumTmp[36][4] , \u_div/SumTmp[37][1] , \u_div/SumTmp[37][2] ,
         \u_div/SumTmp[37][3] , \u_div/SumTmp[37][4] , \u_div/SumTmp[38][1] ,
         \u_div/SumTmp[38][2] , \u_div/SumTmp[38][3] , \u_div/SumTmp[38][4] ,
         \u_div/SumTmp[39][1] , \u_div/SumTmp[39][2] , \u_div/SumTmp[39][3] ,
         \u_div/SumTmp[39][4] , \u_div/SumTmp[40][1] , \u_div/SumTmp[40][2] ,
         \u_div/SumTmp[40][3] , \u_div/SumTmp[40][4] , \u_div/SumTmp[41][1] ,
         \u_div/SumTmp[41][2] , \u_div/SumTmp[41][3] , \u_div/SumTmp[41][4] ,
         \u_div/SumTmp[42][1] , \u_div/SumTmp[42][2] , \u_div/SumTmp[42][3] ,
         \u_div/SumTmp[42][4] , \u_div/SumTmp[43][1] , \u_div/SumTmp[43][2] ,
         \u_div/SumTmp[43][3] , \u_div/SumTmp[43][4] , \u_div/SumTmp[44][1] ,
         \u_div/SumTmp[44][2] , \u_div/SumTmp[44][3] , \u_div/SumTmp[44][4] ,
         \u_div/SumTmp[45][1] , \u_div/SumTmp[45][2] , \u_div/SumTmp[45][3] ,
         \u_div/SumTmp[45][4] , \u_div/SumTmp[46][1] , \u_div/SumTmp[46][2] ,
         \u_div/SumTmp[46][3] , \u_div/SumTmp[46][4] , \u_div/SumTmp[47][1] ,
         \u_div/SumTmp[47][2] , \u_div/SumTmp[47][3] , \u_div/SumTmp[47][4] ,
         \u_div/SumTmp[48][1] , \u_div/SumTmp[48][2] , \u_div/SumTmp[48][3] ,
         \u_div/SumTmp[48][4] , \u_div/SumTmp[49][1] , \u_div/SumTmp[49][2] ,
         \u_div/SumTmp[49][3] , \u_div/SumTmp[49][4] , \u_div/SumTmp[50][1] ,
         \u_div/SumTmp[50][2] , \u_div/SumTmp[50][3] , \u_div/SumTmp[50][4] ,
         \u_div/SumTmp[51][1] , \u_div/SumTmp[51][2] , \u_div/SumTmp[51][3] ,
         \u_div/SumTmp[51][4] , \u_div/SumTmp[52][1] , \u_div/SumTmp[52][2] ,
         \u_div/SumTmp[52][3] , \u_div/SumTmp[52][4] , \u_div/SumTmp[53][1] ,
         \u_div/SumTmp[53][2] , \u_div/SumTmp[53][3] , \u_div/SumTmp[53][4] ,
         \u_div/SumTmp[54][1] , \u_div/SumTmp[54][2] , \u_div/SumTmp[54][3] ,
         \u_div/SumTmp[54][4] , \u_div/SumTmp[55][1] , \u_div/SumTmp[55][2] ,
         \u_div/SumTmp[55][3] , \u_div/SumTmp[55][4] , \u_div/SumTmp[56][1] ,
         \u_div/SumTmp[56][2] , \u_div/SumTmp[56][3] , \u_div/SumTmp[56][4] ,
         \u_div/SumTmp[57][1] , \u_div/SumTmp[57][2] , \u_div/SumTmp[57][3] ,
         \u_div/SumTmp[57][4] , \u_div/SumTmp[58][1] , \u_div/SumTmp[58][2] ,
         \u_div/SumTmp[58][3] , \u_div/SumTmp[58][4] , \u_div/SumTmp[59][3] ,
         \u_div/SumTmp[59][4] , \u_div/CryTmp[0][6] , \u_div/CryTmp[1][6] ,
         \u_div/CryTmp[2][6] , \u_div/CryTmp[3][6] , \u_div/CryTmp[4][6] ,
         \u_div/CryTmp[5][6] , \u_div/CryTmp[6][6] , \u_div/CryTmp[7][6] ,
         \u_div/CryTmp[8][6] , \u_div/CryTmp[9][6] , \u_div/CryTmp[10][6] ,
         \u_div/CryTmp[11][6] , \u_div/CryTmp[12][6] , \u_div/CryTmp[13][6] ,
         \u_div/CryTmp[14][6] , \u_div/CryTmp[15][6] , \u_div/CryTmp[16][6] ,
         \u_div/CryTmp[17][6] , \u_div/CryTmp[18][6] , \u_div/CryTmp[19][6] ,
         \u_div/CryTmp[20][6] , \u_div/CryTmp[21][6] , \u_div/CryTmp[22][6] ,
         \u_div/CryTmp[23][6] , \u_div/CryTmp[24][6] , \u_div/CryTmp[25][6] ,
         \u_div/CryTmp[26][6] , \u_div/CryTmp[27][6] , \u_div/CryTmp[28][6] ,
         \u_div/CryTmp[29][6] , \u_div/CryTmp[30][6] , \u_div/CryTmp[31][6] ,
         \u_div/CryTmp[32][6] , \u_div/CryTmp[33][6] , \u_div/CryTmp[34][6] ,
         \u_div/CryTmp[35][6] , \u_div/CryTmp[36][6] , \u_div/CryTmp[37][6] ,
         \u_div/CryTmp[38][6] , \u_div/CryTmp[39][6] , \u_div/CryTmp[40][6] ,
         \u_div/CryTmp[41][6] , \u_div/CryTmp[42][6] , \u_div/CryTmp[43][6] ,
         \u_div/CryTmp[44][6] , \u_div/CryTmp[45][6] , \u_div/CryTmp[46][6] ,
         \u_div/CryTmp[47][6] , \u_div/CryTmp[48][6] , \u_div/CryTmp[49][6] ,
         \u_div/CryTmp[50][6] , \u_div/CryTmp[51][6] , \u_div/CryTmp[52][6] ,
         \u_div/CryTmp[53][6] , \u_div/CryTmp[54][6] , \u_div/CryTmp[55][6] ,
         \u_div/CryTmp[56][6] , \u_div/CryTmp[57][6] , \u_div/CryTmp[58][6] ,
         \u_div/CryTmp[59][6] , \u_div/PartRem[1][2] , \u_div/PartRem[1][3] ,
         \u_div/PartRem[1][4] , \u_div/PartRem[1][5] , \u_div/PartRem[2][2] ,
         \u_div/PartRem[2][3] , \u_div/PartRem[2][4] , \u_div/PartRem[2][5] ,
         \u_div/PartRem[3][0] , \u_div/PartRem[3][2] , \u_div/PartRem[3][3] ,
         \u_div/PartRem[3][4] , \u_div/PartRem[3][5] , \u_div/PartRem[4][0] ,
         \u_div/PartRem[4][2] , \u_div/PartRem[4][3] , \u_div/PartRem[4][4] ,
         \u_div/PartRem[4][5] , \u_div/PartRem[5][0] , \u_div/PartRem[5][2] ,
         \u_div/PartRem[5][3] , \u_div/PartRem[5][4] , \u_div/PartRem[5][5] ,
         \u_div/PartRem[6][0] , \u_div/PartRem[6][2] , \u_div/PartRem[6][3] ,
         \u_div/PartRem[6][4] , \u_div/PartRem[6][5] , \u_div/PartRem[7][0] ,
         \u_div/PartRem[7][2] , \u_div/PartRem[7][3] , \u_div/PartRem[7][4] ,
         \u_div/PartRem[7][5] , \u_div/PartRem[8][0] , \u_div/PartRem[8][2] ,
         \u_div/PartRem[8][3] , \u_div/PartRem[8][4] , \u_div/PartRem[8][5] ,
         \u_div/PartRem[9][0] , \u_div/PartRem[9][2] , \u_div/PartRem[9][3] ,
         \u_div/PartRem[9][4] , \u_div/PartRem[9][5] , \u_div/PartRem[10][0] ,
         \u_div/PartRem[10][2] , \u_div/PartRem[10][3] ,
         \u_div/PartRem[10][4] , \u_div/PartRem[10][5] ,
         \u_div/PartRem[11][0] , \u_div/PartRem[11][2] ,
         \u_div/PartRem[11][3] , \u_div/PartRem[11][4] ,
         \u_div/PartRem[11][5] , \u_div/PartRem[12][0] ,
         \u_div/PartRem[12][2] , \u_div/PartRem[12][3] ,
         \u_div/PartRem[12][4] , \u_div/PartRem[12][5] ,
         \u_div/PartRem[13][0] , \u_div/PartRem[13][2] ,
         \u_div/PartRem[13][3] , \u_div/PartRem[13][4] ,
         \u_div/PartRem[13][5] , \u_div/PartRem[14][0] ,
         \u_div/PartRem[14][2] , \u_div/PartRem[14][3] ,
         \u_div/PartRem[14][4] , \u_div/PartRem[14][5] ,
         \u_div/PartRem[15][0] , \u_div/PartRem[15][2] ,
         \u_div/PartRem[15][3] , \u_div/PartRem[15][4] ,
         \u_div/PartRem[15][5] , \u_div/PartRem[16][0] ,
         \u_div/PartRem[16][2] , \u_div/PartRem[16][3] ,
         \u_div/PartRem[16][4] , \u_div/PartRem[16][5] ,
         \u_div/PartRem[17][0] , \u_div/PartRem[17][2] ,
         \u_div/PartRem[17][3] , \u_div/PartRem[17][4] ,
         \u_div/PartRem[17][5] , \u_div/PartRem[18][0] ,
         \u_div/PartRem[18][2] , \u_div/PartRem[18][3] ,
         \u_div/PartRem[18][4] , \u_div/PartRem[18][5] ,
         \u_div/PartRem[19][0] , \u_div/PartRem[19][2] ,
         \u_div/PartRem[19][3] , \u_div/PartRem[19][4] ,
         \u_div/PartRem[19][5] , \u_div/PartRem[20][0] ,
         \u_div/PartRem[20][2] , \u_div/PartRem[20][3] ,
         \u_div/PartRem[20][4] , \u_div/PartRem[20][5] ,
         \u_div/PartRem[21][0] , \u_div/PartRem[21][2] ,
         \u_div/PartRem[21][3] , \u_div/PartRem[21][4] ,
         \u_div/PartRem[21][5] , \u_div/PartRem[22][0] ,
         \u_div/PartRem[22][2] , \u_div/PartRem[22][3] ,
         \u_div/PartRem[22][4] , \u_div/PartRem[22][5] ,
         \u_div/PartRem[23][0] , \u_div/PartRem[23][2] ,
         \u_div/PartRem[23][3] , \u_div/PartRem[23][4] ,
         \u_div/PartRem[23][5] , \u_div/PartRem[24][0] ,
         \u_div/PartRem[24][2] , \u_div/PartRem[24][3] ,
         \u_div/PartRem[24][4] , \u_div/PartRem[24][5] ,
         \u_div/PartRem[25][0] , \u_div/PartRem[25][2] ,
         \u_div/PartRem[25][3] , \u_div/PartRem[25][4] ,
         \u_div/PartRem[25][5] , \u_div/PartRem[26][0] ,
         \u_div/PartRem[26][2] , \u_div/PartRem[26][3] ,
         \u_div/PartRem[26][4] , \u_div/PartRem[26][5] ,
         \u_div/PartRem[27][0] , \u_div/PartRem[27][2] ,
         \u_div/PartRem[27][3] , \u_div/PartRem[27][4] ,
         \u_div/PartRem[27][5] , \u_div/PartRem[28][0] ,
         \u_div/PartRem[28][2] , \u_div/PartRem[28][3] ,
         \u_div/PartRem[28][4] , \u_div/PartRem[28][5] ,
         \u_div/PartRem[29][0] , \u_div/PartRem[29][2] ,
         \u_div/PartRem[29][3] , \u_div/PartRem[29][4] ,
         \u_div/PartRem[29][5] , \u_div/PartRem[30][0] ,
         \u_div/PartRem[30][2] , \u_div/PartRem[30][3] ,
         \u_div/PartRem[30][4] , \u_div/PartRem[30][5] ,
         \u_div/PartRem[31][0] , \u_div/PartRem[31][2] ,
         \u_div/PartRem[31][3] , \u_div/PartRem[31][4] ,
         \u_div/PartRem[31][5] , \u_div/PartRem[32][0] ,
         \u_div/PartRem[32][2] , \u_div/PartRem[32][3] ,
         \u_div/PartRem[32][4] , \u_div/PartRem[32][5] ,
         \u_div/PartRem[33][0] , \u_div/PartRem[33][2] ,
         \u_div/PartRem[33][3] , \u_div/PartRem[33][4] ,
         \u_div/PartRem[33][5] , \u_div/PartRem[34][0] ,
         \u_div/PartRem[34][2] , \u_div/PartRem[34][3] ,
         \u_div/PartRem[34][4] , \u_div/PartRem[34][5] ,
         \u_div/PartRem[35][0] , \u_div/PartRem[35][2] ,
         \u_div/PartRem[35][3] , \u_div/PartRem[35][4] ,
         \u_div/PartRem[35][5] , \u_div/PartRem[36][0] ,
         \u_div/PartRem[36][2] , \u_div/PartRem[36][3] ,
         \u_div/PartRem[36][4] , \u_div/PartRem[36][5] ,
         \u_div/PartRem[37][0] , \u_div/PartRem[37][2] ,
         \u_div/PartRem[37][3] , \u_div/PartRem[37][4] ,
         \u_div/PartRem[37][5] , \u_div/PartRem[38][0] ,
         \u_div/PartRem[38][2] , \u_div/PartRem[38][3] ,
         \u_div/PartRem[38][4] , \u_div/PartRem[38][5] ,
         \u_div/PartRem[39][0] , \u_div/PartRem[39][2] ,
         \u_div/PartRem[39][3] , \u_div/PartRem[39][4] ,
         \u_div/PartRem[39][5] , \u_div/PartRem[40][0] ,
         \u_div/PartRem[40][2] , \u_div/PartRem[40][3] ,
         \u_div/PartRem[40][4] , \u_div/PartRem[40][5] ,
         \u_div/PartRem[41][0] , \u_div/PartRem[41][2] ,
         \u_div/PartRem[41][3] , \u_div/PartRem[41][4] ,
         \u_div/PartRem[41][5] , \u_div/PartRem[42][0] ,
         \u_div/PartRem[42][2] , \u_div/PartRem[42][3] ,
         \u_div/PartRem[42][4] , \u_div/PartRem[42][5] ,
         \u_div/PartRem[43][0] , \u_div/PartRem[43][2] ,
         \u_div/PartRem[43][3] , \u_div/PartRem[43][4] ,
         \u_div/PartRem[43][5] , \u_div/PartRem[44][0] ,
         \u_div/PartRem[44][2] , \u_div/PartRem[44][3] ,
         \u_div/PartRem[44][4] , \u_div/PartRem[44][5] ,
         \u_div/PartRem[45][0] , \u_div/PartRem[45][2] ,
         \u_div/PartRem[45][3] , \u_div/PartRem[45][4] ,
         \u_div/PartRem[45][5] , \u_div/PartRem[46][0] ,
         \u_div/PartRem[46][2] , \u_div/PartRem[46][3] ,
         \u_div/PartRem[46][4] , \u_div/PartRem[46][5] ,
         \u_div/PartRem[47][0] , \u_div/PartRem[47][2] ,
         \u_div/PartRem[47][3] , \u_div/PartRem[47][4] ,
         \u_div/PartRem[47][5] , \u_div/PartRem[48][0] ,
         \u_div/PartRem[48][2] , \u_div/PartRem[48][3] ,
         \u_div/PartRem[48][4] , \u_div/PartRem[48][5] ,
         \u_div/PartRem[49][0] , \u_div/PartRem[49][2] ,
         \u_div/PartRem[49][3] , \u_div/PartRem[49][4] ,
         \u_div/PartRem[49][5] , \u_div/PartRem[50][0] ,
         \u_div/PartRem[50][2] , \u_div/PartRem[50][3] ,
         \u_div/PartRem[50][4] , \u_div/PartRem[50][5] ,
         \u_div/PartRem[51][0] , \u_div/PartRem[51][2] ,
         \u_div/PartRem[51][3] , \u_div/PartRem[51][4] ,
         \u_div/PartRem[51][5] , \u_div/PartRem[52][0] ,
         \u_div/PartRem[52][2] , \u_div/PartRem[52][3] ,
         \u_div/PartRem[52][4] , \u_div/PartRem[52][5] ,
         \u_div/PartRem[53][0] , \u_div/PartRem[53][2] ,
         \u_div/PartRem[53][3] , \u_div/PartRem[53][4] ,
         \u_div/PartRem[53][5] , \u_div/PartRem[54][0] ,
         \u_div/PartRem[54][2] , \u_div/PartRem[54][3] ,
         \u_div/PartRem[54][4] , \u_div/PartRem[54][5] ,
         \u_div/PartRem[55][0] , \u_div/PartRem[55][2] ,
         \u_div/PartRem[55][3] , \u_div/PartRem[55][4] ,
         \u_div/PartRem[55][5] , \u_div/PartRem[56][0] ,
         \u_div/PartRem[56][2] , \u_div/PartRem[56][3] ,
         \u_div/PartRem[56][4] , \u_div/PartRem[56][5] ,
         \u_div/PartRem[57][0] , \u_div/PartRem[57][2] ,
         \u_div/PartRem[57][3] , \u_div/PartRem[57][4] ,
         \u_div/PartRem[57][5] , \u_div/PartRem[58][0] ,
         \u_div/PartRem[58][2] , \u_div/PartRem[58][3] ,
         \u_div/PartRem[58][4] , \u_div/PartRem[58][5] ,
         \u_div/PartRem[59][0] , \u_div/PartRem[59][2] ,
         \u_div/PartRem[59][3] , \u_div/PartRem[59][4] ,
         \u_div/PartRem[59][5] , \u_div/PartRem[60][0] ,
         \u_div/PartRem[61][0] , \u_div/PartRem[62][0] ,
         \u_div/PartRem[63][0] , \u_div/PartRem[64][0] ,
         \u_div/u_add_PartRem_2_1/n3 , \u_div/u_add_PartRem_2_1/n2 ,
         \u_div/u_add_PartRem_2_2/n3 , \u_div/u_add_PartRem_2_2/n2 ,
         \u_div/u_add_PartRem_2_3/n3 , \u_div/u_add_PartRem_2_3/n2 ,
         \u_div/u_add_PartRem_2_4/n3 , \u_div/u_add_PartRem_2_4/n2 ,
         \u_div/u_add_PartRem_2_5/n3 , \u_div/u_add_PartRem_2_5/n2 ,
         \u_div/u_add_PartRem_2_6/n3 , \u_div/u_add_PartRem_2_6/n2 ,
         \u_div/u_add_PartRem_2_7/n3 , \u_div/u_add_PartRem_2_7/n2 ,
         \u_div/u_add_PartRem_2_8/n3 , \u_div/u_add_PartRem_2_8/n2 ,
         \u_div/u_add_PartRem_2_9/n3 , \u_div/u_add_PartRem_2_9/n2 ,
         \u_div/u_add_PartRem_2_10/n3 , \u_div/u_add_PartRem_2_10/n2 ,
         \u_div/u_add_PartRem_2_11/n3 , \u_div/u_add_PartRem_2_11/n2 ,
         \u_div/u_add_PartRem_2_12/n3 , \u_div/u_add_PartRem_2_12/n2 ,
         \u_div/u_add_PartRem_2_13/n3 , \u_div/u_add_PartRem_2_13/n2 ,
         \u_div/u_add_PartRem_2_14/n3 , \u_div/u_add_PartRem_2_14/n2 ,
         \u_div/u_add_PartRem_2_15/n3 , \u_div/u_add_PartRem_2_15/n2 ,
         \u_div/u_add_PartRem_2_16/n3 , \u_div/u_add_PartRem_2_16/n2 ,
         \u_div/u_add_PartRem_2_17/n3 , \u_div/u_add_PartRem_2_17/n2 ,
         \u_div/u_add_PartRem_2_18/n3 , \u_div/u_add_PartRem_2_18/n2 ,
         \u_div/u_add_PartRem_2_19/n3 , \u_div/u_add_PartRem_2_19/n2 ,
         \u_div/u_add_PartRem_2_20/n3 , \u_div/u_add_PartRem_2_20/n2 ,
         \u_div/u_add_PartRem_2_21/n3 , \u_div/u_add_PartRem_2_21/n2 ,
         \u_div/u_add_PartRem_2_22/n3 , \u_div/u_add_PartRem_2_22/n2 ,
         \u_div/u_add_PartRem_2_23/n3 , \u_div/u_add_PartRem_2_23/n2 ,
         \u_div/u_add_PartRem_2_24/n3 , \u_div/u_add_PartRem_2_24/n2 ,
         \u_div/u_add_PartRem_2_25/n3 , \u_div/u_add_PartRem_2_25/n2 ,
         \u_div/u_add_PartRem_2_26/n3 , \u_div/u_add_PartRem_2_26/n2 ,
         \u_div/u_add_PartRem_2_27/n3 , \u_div/u_add_PartRem_2_27/n2 ,
         \u_div/u_add_PartRem_2_28/n3 , \u_div/u_add_PartRem_2_28/n2 ,
         \u_div/u_add_PartRem_2_29/n3 , \u_div/u_add_PartRem_2_29/n2 ,
         \u_div/u_add_PartRem_2_30/n3 , \u_div/u_add_PartRem_2_30/n2 ,
         \u_div/u_add_PartRem_2_31/n3 , \u_div/u_add_PartRem_2_31/n2 ,
         \u_div/u_add_PartRem_2_32/n3 , \u_div/u_add_PartRem_2_32/n2 ,
         \u_div/u_add_PartRem_2_33/n3 , \u_div/u_add_PartRem_2_33/n2 ,
         \u_div/u_add_PartRem_2_34/n3 , \u_div/u_add_PartRem_2_34/n2 ,
         \u_div/u_add_PartRem_2_35/n3 , \u_div/u_add_PartRem_2_35/n2 ,
         \u_div/u_add_PartRem_2_36/n3 , \u_div/u_add_PartRem_2_36/n2 ,
         \u_div/u_add_PartRem_2_37/n3 , \u_div/u_add_PartRem_2_37/n2 ,
         \u_div/u_add_PartRem_2_38/n3 , \u_div/u_add_PartRem_2_38/n2 ,
         \u_div/u_add_PartRem_2_39/n3 , \u_div/u_add_PartRem_2_39/n2 ,
         \u_div/u_add_PartRem_2_40/n3 , \u_div/u_add_PartRem_2_40/n2 ,
         \u_div/u_add_PartRem_2_41/n3 , \u_div/u_add_PartRem_2_41/n2 ,
         \u_div/u_add_PartRem_2_42/n3 , \u_div/u_add_PartRem_2_42/n2 ,
         \u_div/u_add_PartRem_2_43/n3 , \u_div/u_add_PartRem_2_43/n2 ,
         \u_div/u_add_PartRem_2_44/n3 , \u_div/u_add_PartRem_2_44/n2 ,
         \u_div/u_add_PartRem_2_45/n3 , \u_div/u_add_PartRem_2_45/n2 ,
         \u_div/u_add_PartRem_2_46/n3 , \u_div/u_add_PartRem_2_46/n2 ,
         \u_div/u_add_PartRem_2_47/n3 , \u_div/u_add_PartRem_2_47/n2 ,
         \u_div/u_add_PartRem_2_48/n3 , \u_div/u_add_PartRem_2_48/n2 ,
         \u_div/u_add_PartRem_2_49/n3 , \u_div/u_add_PartRem_2_49/n2 ,
         \u_div/u_add_PartRem_2_50/n3 , \u_div/u_add_PartRem_2_50/n2 ,
         \u_div/u_add_PartRem_2_51/n3 , \u_div/u_add_PartRem_2_51/n2 ,
         \u_div/u_add_PartRem_2_52/n3 , \u_div/u_add_PartRem_2_52/n2 ,
         \u_div/u_add_PartRem_2_53/n3 , \u_div/u_add_PartRem_2_53/n2 ,
         \u_div/u_add_PartRem_2_54/n3 , \u_div/u_add_PartRem_2_54/n2 ,
         \u_div/u_add_PartRem_2_55/n3 , \u_div/u_add_PartRem_2_55/n2 ,
         \u_div/u_add_PartRem_2_56/n3 , \u_div/u_add_PartRem_2_56/n2 ,
         \u_div/u_add_PartRem_2_57/n3 , \u_div/u_add_PartRem_2_57/n2 ,
         \u_div/u_add_PartRem_2_58/n3 , \u_div/u_add_PartRem_2_58/n2 , n1, n2,
         n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign \u_div/QInv[63]  = a[63];

  GSIM_DW01_absval_5 \u_div/u_absval_AAbs  ( .A({n2, a[62:0]}), .ABSVAL({
        \u_div/PartRem[64][0] , \u_div/PartRem[63][0] , \u_div/PartRem[62][0] , 
        \u_div/PartRem[61][0] , \u_div/PartRem[60][0] , \u_div/PartRem[59][0] , 
        \u_div/PartRem[58][0] , \u_div/PartRem[57][0] , \u_div/PartRem[56][0] , 
        \u_div/PartRem[55][0] , \u_div/PartRem[54][0] , \u_div/PartRem[53][0] , 
        \u_div/PartRem[52][0] , \u_div/PartRem[51][0] , \u_div/PartRem[50][0] , 
        \u_div/PartRem[49][0] , \u_div/PartRem[48][0] , \u_div/PartRem[47][0] , 
        \u_div/PartRem[46][0] , \u_div/PartRem[45][0] , \u_div/PartRem[44][0] , 
        \u_div/PartRem[43][0] , \u_div/PartRem[42][0] , \u_div/PartRem[41][0] , 
        \u_div/PartRem[40][0] , \u_div/PartRem[39][0] , \u_div/PartRem[38][0] , 
        \u_div/PartRem[37][0] , \u_div/PartRem[36][0] , \u_div/PartRem[35][0] , 
        \u_div/PartRem[34][0] , \u_div/PartRem[33][0] , \u_div/PartRem[32][0] , 
        \u_div/PartRem[31][0] , \u_div/PartRem[30][0] , \u_div/PartRem[29][0] , 
        \u_div/PartRem[28][0] , \u_div/PartRem[27][0] , \u_div/PartRem[26][0] , 
        \u_div/PartRem[25][0] , \u_div/PartRem[24][0] , \u_div/PartRem[23][0] , 
        \u_div/PartRem[22][0] , \u_div/PartRem[21][0] , \u_div/PartRem[20][0] , 
        \u_div/PartRem[19][0] , \u_div/PartRem[18][0] , \u_div/PartRem[17][0] , 
        \u_div/PartRem[16][0] , \u_div/PartRem[15][0] , \u_div/PartRem[14][0] , 
        \u_div/PartRem[13][0] , \u_div/PartRem[12][0] , \u_div/PartRem[11][0] , 
        \u_div/PartRem[10][0] , \u_div/PartRem[9][0] , \u_div/PartRem[8][0] , 
        \u_div/PartRem[7][0] , \u_div/PartRem[6][0] , \u_div/PartRem[5][0] , 
        \u_div/PartRem[4][0] , \u_div/PartRem[3][0] , SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1}) );
  GSIM_DW_inc_5 \u_div/u_inc_QInc  ( .carry_in(n4), .a({n2, n2, n2, n3, 
        \u_div/QInv[59] , \u_div/QInv[58] , \u_div/QInv[57] , \u_div/QInv[56] , 
        \u_div/QInv[55] , \u_div/QInv[54] , \u_div/QInv[53] , \u_div/QInv[52] , 
        \u_div/QInv[51] , \u_div/QInv[50] , \u_div/QInv[49] , \u_div/QInv[48] , 
        \u_div/QInv[47] , \u_div/QInv[46] , \u_div/QInv[45] , \u_div/QInv[44] , 
        \u_div/QInv[43] , \u_div/QInv[42] , \u_div/QInv[41] , \u_div/QInv[40] , 
        \u_div/QInv[39] , \u_div/QInv[38] , \u_div/QInv[37] , \u_div/QInv[36] , 
        \u_div/QInv[35] , \u_div/QInv[34] , \u_div/QInv[33] , \u_div/QInv[32] , 
        \u_div/QInv[31] , \u_div/QInv[30] , \u_div/QInv[29] , \u_div/QInv[28] , 
        \u_div/QInv[27] , \u_div/QInv[26] , \u_div/QInv[25] , \u_div/QInv[24] , 
        \u_div/QInv[23] , \u_div/QInv[22] , \u_div/QInv[21] , \u_div/QInv[20] , 
        \u_div/QInv[19] , \u_div/QInv[18] , \u_div/QInv[17] , \u_div/QInv[16] , 
        \u_div/QInv[15] , \u_div/QInv[14] , \u_div/QInv[13] , \u_div/QInv[12] , 
        \u_div/QInv[11] , \u_div/QInv[10] , \u_div/QInv[9] , \u_div/QInv[8] , 
        \u_div/QInv[7] , \u_div/QInv[6] , \u_div/QInv[5] , \u_div/QInv[4] , 
        \u_div/QInv[3] , \u_div/QInv[2] , \u_div/QInv[1] , \u_div/QInv[0] }), 
        .sum(quotient) );
  ADDHXL \u_div/u_add_PartRem_2_6/U3  ( .A(\u_div/PartRem[7][4] ), .B(
        \u_div/u_add_PartRem_2_6/n3 ), .CO(\u_div/u_add_PartRem_2_6/n2 ), .S(
        \u_div/SumTmp[6][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_11/U3  ( .A(\u_div/PartRem[12][4] ), .B(
        \u_div/u_add_PartRem_2_11/n3 ), .CO(\u_div/u_add_PartRem_2_11/n2 ), 
        .S(\u_div/SumTmp[11][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_16/U3  ( .A(\u_div/PartRem[17][4] ), .B(
        \u_div/u_add_PartRem_2_16/n3 ), .CO(\u_div/u_add_PartRem_2_16/n2 ), 
        .S(\u_div/SumTmp[16][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_21/U3  ( .A(\u_div/PartRem[22][4] ), .B(
        \u_div/u_add_PartRem_2_21/n3 ), .CO(\u_div/u_add_PartRem_2_21/n2 ), 
        .S(\u_div/SumTmp[21][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_26/U3  ( .A(\u_div/PartRem[27][4] ), .B(
        \u_div/u_add_PartRem_2_26/n3 ), .CO(\u_div/u_add_PartRem_2_26/n2 ), 
        .S(\u_div/SumTmp[26][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_31/U3  ( .A(\u_div/PartRem[32][4] ), .B(
        \u_div/u_add_PartRem_2_31/n3 ), .CO(\u_div/u_add_PartRem_2_31/n2 ), 
        .S(\u_div/SumTmp[31][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_36/U3  ( .A(\u_div/PartRem[37][4] ), .B(
        \u_div/u_add_PartRem_2_36/n3 ), .CO(\u_div/u_add_PartRem_2_36/n2 ), 
        .S(\u_div/SumTmp[36][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_41/U3  ( .A(\u_div/PartRem[42][4] ), .B(
        \u_div/u_add_PartRem_2_41/n3 ), .CO(\u_div/u_add_PartRem_2_41/n2 ), 
        .S(\u_div/SumTmp[41][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_46/U3  ( .A(\u_div/PartRem[47][4] ), .B(
        \u_div/u_add_PartRem_2_46/n3 ), .CO(\u_div/u_add_PartRem_2_46/n2 ), 
        .S(\u_div/SumTmp[46][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_51/U3  ( .A(\u_div/PartRem[52][4] ), .B(
        \u_div/u_add_PartRem_2_51/n3 ), .CO(\u_div/u_add_PartRem_2_51/n2 ), 
        .S(\u_div/SumTmp[51][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_56/U3  ( .A(\u_div/PartRem[57][4] ), .B(
        \u_div/u_add_PartRem_2_56/n3 ), .CO(\u_div/u_add_PartRem_2_56/n2 ), 
        .S(\u_div/SumTmp[56][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_0  ( .A(\u_div/PartRem[5][0] ), .B(
        \u_div/PartRem[5][0] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/SumTmp[3][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_3_1  ( .A(\u_div/SumTmp[3][1] ), .B(
        \u_div/SumTmp[3][1] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_0  ( .A(\u_div/PartRem[6][0] ), .B(
        \u_div/PartRem[6][0] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/SumTmp[4][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_0  ( .A(\u_div/PartRem[7][0] ), .B(
        \u_div/PartRem[7][0] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/SumTmp[5][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_0  ( .A(\u_div/PartRem[8][0] ), .B(
        \u_div/PartRem[8][0] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/SumTmp[6][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_9_0  ( .A(\u_div/PartRem[10][0] ), .B(
        \u_div/PartRem[10][0] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/SumTmp[8][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_0  ( .A(\u_div/PartRem[11][0] ), .B(
        \u_div/PartRem[11][0] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/SumTmp[9][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_0  ( .A(\u_div/PartRem[12][0] ), .B(
        \u_div/PartRem[12][0] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/SumTmp[10][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_0  ( .A(\u_div/PartRem[13][0] ), .B(
        \u_div/PartRem[13][0] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/SumTmp[11][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_0  ( .A(\u_div/PartRem[15][0] ), .B(
        \u_div/PartRem[15][0] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/SumTmp[13][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_0  ( .A(\u_div/PartRem[16][0] ), .B(
        \u_div/PartRem[16][0] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/SumTmp[14][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_0  ( .A(\u_div/PartRem[17][0] ), .B(
        \u_div/PartRem[17][0] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/SumTmp[15][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_0  ( .A(\u_div/PartRem[18][0] ), .B(
        \u_div/PartRem[18][0] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/SumTmp[16][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_0  ( .A(\u_div/PartRem[20][0] ), .B(
        \u_div/PartRem[20][0] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/SumTmp[18][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_0  ( .A(\u_div/PartRem[21][0] ), .B(
        \u_div/PartRem[21][0] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/SumTmp[19][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_0  ( .A(\u_div/PartRem[22][0] ), .B(
        \u_div/PartRem[22][0] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/SumTmp[20][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_0  ( .A(\u_div/PartRem[23][0] ), .B(
        \u_div/PartRem[23][0] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/SumTmp[21][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_0  ( .A(\u_div/PartRem[25][0] ), .B(
        \u_div/PartRem[25][0] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/SumTmp[23][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_0  ( .A(\u_div/PartRem[26][0] ), .B(
        \u_div/PartRem[26][0] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/SumTmp[24][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_0  ( .A(\u_div/PartRem[27][0] ), .B(
        \u_div/PartRem[27][0] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/SumTmp[25][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_0  ( .A(\u_div/PartRem[28][0] ), .B(
        \u_div/PartRem[28][0] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/SumTmp[26][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_0  ( .A(\u_div/PartRem[30][0] ), .B(
        \u_div/PartRem[30][0] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/SumTmp[28][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_0  ( .A(\u_div/PartRem[31][0] ), .B(
        \u_div/PartRem[31][0] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/SumTmp[29][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_0  ( .A(\u_div/PartRem[32][0] ), .B(
        \u_div/PartRem[32][0] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/SumTmp[30][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_0  ( .A(\u_div/PartRem[33][0] ), .B(
        \u_div/PartRem[33][0] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/SumTmp[31][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_0  ( .A(\u_div/PartRem[35][0] ), .B(
        \u_div/PartRem[35][0] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/SumTmp[33][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_0  ( .A(\u_div/PartRem[36][0] ), .B(
        \u_div/PartRem[36][0] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/SumTmp[34][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_0  ( .A(\u_div/PartRem[37][0] ), .B(
        \u_div/PartRem[37][0] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/SumTmp[35][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_0  ( .A(\u_div/PartRem[38][0] ), .B(
        \u_div/PartRem[38][0] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/SumTmp[36][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_0  ( .A(\u_div/PartRem[40][0] ), .B(
        \u_div/PartRem[40][0] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/SumTmp[38][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_0  ( .A(\u_div/PartRem[41][0] ), .B(
        \u_div/PartRem[41][0] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/SumTmp[39][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_0  ( .A(\u_div/PartRem[42][0] ), .B(
        \u_div/PartRem[42][0] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/SumTmp[40][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_0  ( .A(\u_div/PartRem[43][0] ), .B(
        \u_div/PartRem[43][0] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/SumTmp[41][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_0  ( .A(\u_div/PartRem[45][0] ), .B(
        \u_div/PartRem[45][0] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/SumTmp[43][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_0  ( .A(\u_div/PartRem[46][0] ), .B(
        \u_div/PartRem[46][0] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/SumTmp[44][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_0  ( .A(\u_div/PartRem[47][0] ), .B(
        \u_div/PartRem[47][0] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/SumTmp[45][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_0  ( .A(\u_div/PartRem[48][0] ), .B(
        \u_div/PartRem[48][0] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/SumTmp[46][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_0  ( .A(\u_div/PartRem[50][0] ), .B(
        \u_div/PartRem[50][0] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/SumTmp[48][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_0  ( .A(\u_div/PartRem[51][0] ), .B(
        \u_div/PartRem[51][0] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/SumTmp[49][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_0  ( .A(\u_div/PartRem[52][0] ), .B(
        \u_div/PartRem[52][0] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/SumTmp[50][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_0  ( .A(\u_div/PartRem[53][0] ), .B(
        \u_div/PartRem[53][0] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/SumTmp[51][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_0  ( .A(\u_div/PartRem[55][0] ), .B(
        \u_div/PartRem[55][0] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/SumTmp[53][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_0  ( .A(\u_div/PartRem[56][0] ), .B(
        \u_div/PartRem[56][0] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/SumTmp[54][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_0  ( .A(\u_div/PartRem[57][0] ), .B(
        \u_div/PartRem[57][0] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/SumTmp[55][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_0  ( .A(\u_div/PartRem[58][0] ), .B(
        \u_div/PartRem[58][0] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/SumTmp[56][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_0  ( .A(\u_div/PartRem[60][0] ), .B(
        \u_div/PartRem[60][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/SumTmp[58][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_8_0  ( .A(\u_div/PartRem[9][0] ), .B(
        \u_div/PartRem[9][0] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/SumTmp[7][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_0  ( .A(\u_div/PartRem[19][0] ), .B(
        \u_div/PartRem[19][0] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/SumTmp[17][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_0  ( .A(\u_div/PartRem[29][0] ), .B(
        \u_div/PartRem[29][0] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/SumTmp[27][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_0  ( .A(\u_div/PartRem[34][0] ), .B(
        \u_div/PartRem[34][0] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/SumTmp[32][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_0  ( .A(\u_div/PartRem[39][0] ), .B(
        \u_div/PartRem[39][0] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/SumTmp[37][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_0  ( .A(\u_div/PartRem[44][0] ), .B(
        \u_div/PartRem[44][0] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/SumTmp[42][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_0  ( .A(\u_div/PartRem[49][0] ), .B(
        \u_div/PartRem[49][0] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/SumTmp[47][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_0  ( .A(\u_div/PartRem[54][0] ), .B(
        \u_div/PartRem[54][0] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/SumTmp[52][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_0  ( .A(\u_div/PartRem[59][0] ), .B(
        \u_div/PartRem[59][0] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/SumTmp[57][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_0  ( .A(\u_div/PartRem[14][0] ), .B(
        \u_div/PartRem[14][0] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/SumTmp[12][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_0  ( .A(\u_div/PartRem[24][0] ), .B(
        \u_div/PartRem[24][0] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/SumTmp[22][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_2_1  ( .A(\u_div/SumTmp[2][1] ), .B(
        \u_div/SumTmp[2][1] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_1_1  ( .A(\u_div/SumTmp[1][1] ), .B(
        \u_div/SumTmp[1][1] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_3  ( .A(\u_div/PartRem[5][3] ), .B(
        \u_div/SumTmp[4][3] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_3  ( .A(\u_div/PartRem[6][3] ), .B(
        \u_div/SumTmp[5][3] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_3  ( .A(\u_div/PartRem[7][3] ), .B(
        \u_div/SumTmp[6][3] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_3  ( .A(\u_div/PartRem[8][3] ), .B(
        \u_div/SumTmp[7][3] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_8_3  ( .A(\u_div/PartRem[9][3] ), .B(
        \u_div/SumTmp[8][3] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_9_3  ( .A(\u_div/PartRem[10][3] ), .B(
        \u_div/SumTmp[9][3] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_3  ( .A(\u_div/PartRem[11][3] ), .B(
        \u_div/SumTmp[10][3] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_3  ( .A(\u_div/PartRem[12][3] ), .B(
        \u_div/SumTmp[11][3] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_3  ( .A(\u_div/PartRem[13][3] ), .B(
        \u_div/SumTmp[12][3] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_3  ( .A(\u_div/PartRem[14][3] ), .B(
        \u_div/SumTmp[13][3] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_3  ( .A(\u_div/PartRem[15][3] ), .B(
        \u_div/SumTmp[14][3] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_3  ( .A(\u_div/PartRem[16][3] ), .B(
        \u_div/SumTmp[15][3] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_3  ( .A(\u_div/PartRem[17][3] ), .B(
        \u_div/SumTmp[16][3] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_3  ( .A(\u_div/PartRem[18][3] ), .B(
        \u_div/SumTmp[17][3] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_3  ( .A(\u_div/PartRem[19][3] ), .B(
        \u_div/SumTmp[18][3] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_3  ( .A(\u_div/PartRem[20][3] ), .B(
        \u_div/SumTmp[19][3] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_3  ( .A(\u_div/PartRem[21][3] ), .B(
        \u_div/SumTmp[20][3] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_3  ( .A(\u_div/PartRem[22][3] ), .B(
        \u_div/SumTmp[21][3] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_3  ( .A(\u_div/PartRem[23][3] ), .B(
        \u_div/SumTmp[22][3] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_3  ( .A(\u_div/PartRem[24][3] ), .B(
        \u_div/SumTmp[23][3] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_3  ( .A(\u_div/PartRem[25][3] ), .B(
        \u_div/SumTmp[24][3] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_3  ( .A(\u_div/PartRem[26][3] ), .B(
        \u_div/SumTmp[25][3] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_3  ( .A(\u_div/PartRem[27][3] ), .B(
        \u_div/SumTmp[26][3] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_3  ( .A(\u_div/PartRem[28][3] ), .B(
        \u_div/SumTmp[27][3] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_3  ( .A(\u_div/PartRem[29][3] ), .B(
        \u_div/SumTmp[28][3] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_3  ( .A(\u_div/PartRem[30][3] ), .B(
        \u_div/SumTmp[29][3] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_3  ( .A(\u_div/PartRem[31][3] ), .B(
        \u_div/SumTmp[30][3] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_3  ( .A(\u_div/PartRem[32][3] ), .B(
        \u_div/SumTmp[31][3] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_3  ( .A(\u_div/PartRem[33][3] ), .B(
        \u_div/SumTmp[32][3] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_3  ( .A(\u_div/PartRem[34][3] ), .B(
        \u_div/SumTmp[33][3] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_3  ( .A(\u_div/PartRem[35][3] ), .B(
        \u_div/SumTmp[34][3] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_3  ( .A(\u_div/PartRem[36][3] ), .B(
        \u_div/SumTmp[35][3] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_3  ( .A(\u_div/PartRem[37][3] ), .B(
        \u_div/SumTmp[36][3] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_3  ( .A(\u_div/PartRem[38][3] ), .B(
        \u_div/SumTmp[37][3] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_3  ( .A(\u_div/PartRem[39][3] ), .B(
        \u_div/SumTmp[38][3] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_3  ( .A(\u_div/PartRem[40][3] ), .B(
        \u_div/SumTmp[39][3] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_3  ( .A(\u_div/PartRem[41][3] ), .B(
        \u_div/SumTmp[40][3] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_3  ( .A(\u_div/PartRem[42][3] ), .B(
        \u_div/SumTmp[41][3] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_3  ( .A(\u_div/PartRem[43][3] ), .B(
        \u_div/SumTmp[42][3] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_3  ( .A(\u_div/PartRem[44][3] ), .B(
        \u_div/SumTmp[43][3] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_3  ( .A(\u_div/PartRem[45][3] ), .B(
        \u_div/SumTmp[44][3] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_3  ( .A(\u_div/PartRem[46][3] ), .B(
        \u_div/SumTmp[45][3] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_3  ( .A(\u_div/PartRem[47][3] ), .B(
        \u_div/SumTmp[46][3] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_3  ( .A(\u_div/PartRem[48][3] ), .B(
        \u_div/SumTmp[47][3] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_3  ( .A(\u_div/PartRem[49][3] ), .B(
        \u_div/SumTmp[48][3] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_3  ( .A(\u_div/PartRem[50][3] ), .B(
        \u_div/SumTmp[49][3] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_3  ( .A(\u_div/PartRem[51][3] ), .B(
        \u_div/SumTmp[50][3] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_3  ( .A(\u_div/PartRem[52][3] ), .B(
        \u_div/SumTmp[51][3] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_3  ( .A(\u_div/PartRem[53][3] ), .B(
        \u_div/SumTmp[52][3] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_3  ( .A(\u_div/PartRem[54][3] ), .B(
        \u_div/SumTmp[53][3] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_3  ( .A(\u_div/PartRem[55][3] ), .B(
        \u_div/SumTmp[54][3] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_3  ( .A(\u_div/PartRem[56][3] ), .B(
        \u_div/SumTmp[55][3] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_3  ( .A(\u_div/PartRem[57][3] ), .B(
        \u_div/SumTmp[56][3] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_3  ( .A(\u_div/PartRem[58][3] ), .B(
        \u_div/SumTmp[57][3] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_3  ( .A(\u_div/PartRem[59][3] ), .B(
        \u_div/SumTmp[58][3] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_3  ( .A(\u_div/PartRem[63][0] ), .B(
        \u_div/SumTmp[59][3] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_2_4  ( .A(\u_div/PartRem[3][4] ), .B(
        \u_div/SumTmp[2][4] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_4  ( .A(\u_div/PartRem[64][0] ), .B(
        \u_div/SumTmp[59][4] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_0  ( .A(\u_div/PartRem[3][0] ), .B(
        \u_div/PartRem[3][0] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/SumTmp[1][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_0  ( .A(\u_div/PartRem[4][0] ), .B(
        \u_div/PartRem[4][0] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/SumTmp[2][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_4_1  ( .A(\u_div/SumTmp[4][1] ), .B(
        \u_div/SumTmp[4][1] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_5_1  ( .A(\u_div/SumTmp[5][1] ), .B(
        \u_div/SumTmp[5][1] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_6_1  ( .A(\u_div/SumTmp[6][1] ), .B(
        \u_div/SumTmp[6][1] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_7_1  ( .A(\u_div/SumTmp[7][1] ), .B(
        \u_div/SumTmp[7][1] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_10_1  ( .A(\u_div/SumTmp[10][1] ), .B(
        \u_div/SumTmp[10][1] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_9_1  ( .A(\u_div/SumTmp[9][1] ), .B(
        \u_div/SumTmp[9][1] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_8_1  ( .A(\u_div/SumTmp[8][1] ), .B(
        \u_div/SumTmp[8][1] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_23_1  ( .A(\u_div/SumTmp[23][1] ), .B(
        \u_div/SumTmp[23][1] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_26_1  ( .A(\u_div/SumTmp[26][1] ), .B(
        \u_div/SumTmp[26][1] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_25_1  ( .A(\u_div/SumTmp[25][1] ), .B(
        \u_div/SumTmp[25][1] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_24_1  ( .A(\u_div/SumTmp[24][1] ), .B(
        \u_div/SumTmp[24][1] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_22_1  ( .A(\u_div/SumTmp[22][1] ), .B(
        \u_div/SumTmp[22][1] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_11_1  ( .A(\u_div/SumTmp[11][1] ), .B(
        \u_div/SumTmp[11][1] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_27_1  ( .A(\u_div/SumTmp[27][1] ), .B(
        \u_div/SumTmp[27][1] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_28_1  ( .A(\u_div/SumTmp[28][1] ), .B(
        \u_div/SumTmp[28][1] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_29_1  ( .A(\u_div/SumTmp[29][1] ), .B(
        \u_div/SumTmp[29][1] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_21_1  ( .A(\u_div/SumTmp[21][1] ), .B(
        \u_div/SumTmp[21][1] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_12_1  ( .A(\u_div/SumTmp[12][1] ), .B(
        \u_div/SumTmp[12][1] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_30_1  ( .A(\u_div/SumTmp[30][1] ), .B(
        \u_div/SumTmp[30][1] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_20_1  ( .A(\u_div/SumTmp[20][1] ), .B(
        \u_div/SumTmp[20][1] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_13_1  ( .A(\u_div/SumTmp[13][1] ), .B(
        \u_div/SumTmp[13][1] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_31_1  ( .A(\u_div/SumTmp[31][1] ), .B(
        \u_div/SumTmp[31][1] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_19_1  ( .A(\u_div/SumTmp[19][1] ), .B(
        \u_div/SumTmp[19][1] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_18_1  ( .A(\u_div/SumTmp[18][1] ), .B(
        \u_div/SumTmp[18][1] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_32_1  ( .A(\u_div/SumTmp[32][1] ), .B(
        \u_div/SumTmp[32][1] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_33_1  ( .A(\u_div/SumTmp[33][1] ), .B(
        \u_div/SumTmp[33][1] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_14_1  ( .A(\u_div/SumTmp[14][1] ), .B(
        \u_div/SumTmp[14][1] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_34_1  ( .A(\u_div/SumTmp[34][1] ), .B(
        \u_div/SumTmp[34][1] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_17_1  ( .A(\u_div/SumTmp[17][1] ), .B(
        \u_div/SumTmp[17][1] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_15_1  ( .A(\u_div/SumTmp[15][1] ), .B(
        \u_div/SumTmp[15][1] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_16_1  ( .A(\u_div/SumTmp[16][1] ), .B(
        \u_div/SumTmp[16][1] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_35_1  ( .A(\u_div/SumTmp[35][1] ), .B(
        \u_div/SumTmp[35][1] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_36_1  ( .A(\u_div/SumTmp[36][1] ), .B(
        \u_div/SumTmp[36][1] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_37_1  ( .A(\u_div/SumTmp[37][1] ), .B(
        \u_div/SumTmp[37][1] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_38_1  ( .A(\u_div/SumTmp[38][1] ), .B(
        \u_div/SumTmp[38][1] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_39_1  ( .A(\u_div/SumTmp[39][1] ), .B(
        \u_div/SumTmp[39][1] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_40_1  ( .A(\u_div/SumTmp[40][1] ), .B(
        \u_div/SumTmp[40][1] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_41_1  ( .A(\u_div/SumTmp[41][1] ), .B(
        \u_div/SumTmp[41][1] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_42_1  ( .A(\u_div/SumTmp[42][1] ), .B(
        \u_div/SumTmp[42][1] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_51_1  ( .A(\u_div/SumTmp[51][1] ), .B(
        \u_div/SumTmp[51][1] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_43_1  ( .A(\u_div/SumTmp[43][1] ), .B(
        \u_div/SumTmp[43][1] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_44_1  ( .A(\u_div/SumTmp[44][1] ), .B(
        \u_div/SumTmp[44][1] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_45_1  ( .A(\u_div/SumTmp[45][1] ), .B(
        \u_div/SumTmp[45][1] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_52_1  ( .A(\u_div/SumTmp[52][1] ), .B(
        \u_div/SumTmp[52][1] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_50_1  ( .A(\u_div/SumTmp[50][1] ), .B(
        \u_div/SumTmp[50][1] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_48_1  ( .A(\u_div/SumTmp[48][1] ), .B(
        \u_div/SumTmp[48][1] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_47_1  ( .A(\u_div/SumTmp[47][1] ), .B(
        \u_div/SumTmp[47][1] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_46_1  ( .A(\u_div/SumTmp[46][1] ), .B(
        \u_div/SumTmp[46][1] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_49_1  ( .A(\u_div/SumTmp[49][1] ), .B(
        \u_div/SumTmp[49][1] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_53_1  ( .A(\u_div/SumTmp[53][1] ), .B(
        \u_div/SumTmp[53][1] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_54_1  ( .A(\u_div/SumTmp[54][1] ), .B(
        \u_div/SumTmp[54][1] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_55_1  ( .A(\u_div/SumTmp[55][1] ), .B(
        \u_div/SumTmp[55][1] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_56_1  ( .A(\u_div/SumTmp[56][1] ), .B(
        \u_div/SumTmp[56][1] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_57_1  ( .A(\u_div/SumTmp[57][1] ), .B(
        \u_div/SumTmp[57][1] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_58_1  ( .A(\u_div/SumTmp[58][1] ), .B(
        \u_div/SumTmp[58][1] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_1_3  ( .A(\u_div/PartRem[2][3] ), .B(
        \u_div/SumTmp[1][3] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_3  ( .A(\u_div/PartRem[3][3] ), .B(
        \u_div/SumTmp[2][3] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_3  ( .A(\u_div/PartRem[4][3] ), .B(
        \u_div/SumTmp[3][3] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_1_4  ( .A(\u_div/PartRem[2][4] ), .B(
        \u_div/SumTmp[1][4] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_4  ( .A(\u_div/PartRem[4][4] ), .B(
        \u_div/SumTmp[3][4] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_4  ( .A(\u_div/PartRem[5][4] ), .B(
        \u_div/SumTmp[4][4] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_4  ( .A(\u_div/PartRem[6][4] ), .B(
        \u_div/SumTmp[5][4] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_9_4  ( .A(\u_div/PartRem[10][4] ), .B(
        \u_div/SumTmp[9][4] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_4  ( .A(\u_div/PartRem[7][4] ), .B(
        \u_div/SumTmp[6][4] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_4  ( .A(\u_div/PartRem[26][4] ), .B(
        \u_div/SumTmp[25][4] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_4  ( .A(\u_div/PartRem[23][4] ), .B(
        \u_div/SumTmp[22][4] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_4  ( .A(\u_div/PartRem[11][4] ), .B(
        \u_div/SumTmp[10][4] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_4  ( .A(\u_div/PartRem[8][4] ), .B(
        \u_div/SumTmp[7][4] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_8_4  ( .A(\u_div/PartRem[9][4] ), .B(
        \u_div/SumTmp[8][4] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_4  ( .A(\u_div/PartRem[21][4] ), .B(
        \u_div/SumTmp[20][4] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_4  ( .A(\u_div/PartRem[29][4] ), .B(
        \u_div/SumTmp[28][4] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_4  ( .A(\u_div/PartRem[25][4] ), .B(
        \u_div/SumTmp[24][4] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_4  ( .A(\u_div/PartRem[24][4] ), .B(
        \u_div/SumTmp[23][4] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_4  ( .A(\u_div/PartRem[22][4] ), .B(
        \u_div/SumTmp[21][4] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_4  ( .A(\u_div/PartRem[27][4] ), .B(
        \u_div/SumTmp[26][4] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_4  ( .A(\u_div/PartRem[28][4] ), .B(
        \u_div/SumTmp[27][4] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_4  ( .A(\u_div/PartRem[20][4] ), .B(
        \u_div/SumTmp[19][4] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_4  ( .A(\u_div/PartRem[12][4] ), .B(
        \u_div/SumTmp[11][4] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_4  ( .A(\u_div/PartRem[30][4] ), .B(
        \u_div/SumTmp[29][4] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_4  ( .A(\u_div/PartRem[34][4] ), .B(
        \u_div/SumTmp[33][4] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_4  ( .A(\u_div/PartRem[19][4] ), .B(
        \u_div/SumTmp[18][4] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_4  ( .A(\u_div/PartRem[18][4] ), .B(
        \u_div/SumTmp[17][4] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_4  ( .A(\u_div/PartRem[31][4] ), .B(
        \u_div/SumTmp[30][4] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_4  ( .A(\u_div/PartRem[13][4] ), .B(
        \u_div/SumTmp[12][4] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_4  ( .A(\u_div/PartRem[33][4] ), .B(
        \u_div/SumTmp[32][4] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_4  ( .A(\u_div/PartRem[17][4] ), .B(
        \u_div/SumTmp[16][4] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_4  ( .A(\u_div/PartRem[32][4] ), .B(
        \u_div/SumTmp[31][4] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_4  ( .A(\u_div/PartRem[14][4] ), .B(
        \u_div/SumTmp[13][4] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_4  ( .A(\u_div/PartRem[16][4] ), .B(
        \u_div/SumTmp[15][4] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_4  ( .A(\u_div/PartRem[15][4] ), .B(
        \u_div/SumTmp[14][4] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_4  ( .A(\u_div/PartRem[35][4] ), .B(
        \u_div/SumTmp[34][4] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_4  ( .A(\u_div/PartRem[39][4] ), .B(
        \u_div/SumTmp[38][4] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_4  ( .A(\u_div/PartRem[36][4] ), .B(
        \u_div/SumTmp[35][4] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_4  ( .A(\u_div/PartRem[37][4] ), .B(
        \u_div/SumTmp[36][4] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_4  ( .A(\u_div/PartRem[38][4] ), .B(
        \u_div/SumTmp[37][4] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_4  ( .A(\u_div/PartRem[40][4] ), .B(
        \u_div/SumTmp[39][4] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_4  ( .A(\u_div/PartRem[44][4] ), .B(
        \u_div/SumTmp[43][4] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_4  ( .A(\u_div/PartRem[47][4] ), .B(
        \u_div/SumTmp[46][4] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_4  ( .A(\u_div/PartRem[50][4] ), .B(
        \u_div/SumTmp[49][4] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_4  ( .A(\u_div/PartRem[52][4] ), .B(
        \u_div/SumTmp[51][4] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_4  ( .A(\u_div/PartRem[41][4] ), .B(
        \u_div/SumTmp[40][4] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_4  ( .A(\u_div/PartRem[43][4] ), .B(
        \u_div/SumTmp[42][4] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_4  ( .A(\u_div/PartRem[55][4] ), .B(
        \u_div/SumTmp[54][4] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_4  ( .A(\u_div/PartRem[42][4] ), .B(
        \u_div/SumTmp[41][4] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_4  ( .A(\u_div/PartRem[46][4] ), .B(
        \u_div/SumTmp[45][4] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_4  ( .A(\u_div/PartRem[51][4] ), .B(
        \u_div/SumTmp[50][4] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_4  ( .A(\u_div/PartRem[49][4] ), .B(
        \u_div/SumTmp[48][4] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_4  ( .A(\u_div/PartRem[48][4] ), .B(
        \u_div/SumTmp[47][4] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_4  ( .A(\u_div/PartRem[45][4] ), .B(
        \u_div/SumTmp[44][4] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_4  ( .A(\u_div/PartRem[54][4] ), .B(
        \u_div/SumTmp[53][4] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_4  ( .A(\u_div/PartRem[53][4] ), .B(
        \u_div/SumTmp[52][4] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_4  ( .A(\u_div/PartRem[58][4] ), .B(
        \u_div/SumTmp[57][4] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_4  ( .A(\u_div/PartRem[56][4] ), .B(
        \u_div/SumTmp[55][4] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_4  ( .A(\u_div/PartRem[57][4] ), .B(
        \u_div/SumTmp[56][4] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_4  ( .A(\u_div/PartRem[59][4] ), .B(
        \u_div/SumTmp[58][4] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_59_1  ( .A(\u_div/PartRem[61][0] ), .B(
        \u_div/PartRem[61][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/SumTmp[1][2] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][3] ) );
  OR2X4 U1 ( .A(\u_div/PartRem[17][5] ), .B(\u_div/u_add_PartRem_2_16/n2 ), 
        .Y(\u_div/CryTmp[16][6] ) );
  ADDHXL U2 ( .A(\u_div/PartRem[3][4] ), .B(\u_div/u_add_PartRem_2_2/n3 ), 
        .CO(\u_div/u_add_PartRem_2_2/n2 ), .S(\u_div/SumTmp[2][4] ) );
  INVX3 U3 ( .A(\u_div/QInv[63] ), .Y(n1) );
  OR2X2 U4 ( .A(\u_div/PartRem[12][5] ), .B(\u_div/u_add_PartRem_2_11/n2 ), 
        .Y(\u_div/CryTmp[11][6] ) );
  MXI2X2 U5 ( .A(\u_div/SumTmp[3][2] ), .B(\u_div/PartRem[4][2] ), .S0(
        \u_div/CryTmp[3][6] ), .Y(\u_div/PartRem[3][3] ) );
  OR2X2 U6 ( .A(\u_div/PartRem[22][2] ), .B(\u_div/PartRem[22][3] ), .Y(
        \u_div/u_add_PartRem_2_21/n3 ) );
  OR2X6 U7 ( .A(\u_div/PartRem[3][5] ), .B(\u_div/u_add_PartRem_2_2/n2 ), .Y(
        \u_div/CryTmp[2][6] ) );
  OR2X1 U8 ( .A(\u_div/PartRem[27][2] ), .B(\u_div/PartRem[27][3] ), .Y(
        \u_div/u_add_PartRem_2_26/n3 ) );
  OR2X1 U9 ( .A(\u_div/PartRem[7][2] ), .B(\u_div/PartRem[7][3] ), .Y(
        \u_div/u_add_PartRem_2_6/n3 ) );
  NOR2X6 U10 ( .A(\u_div/PartRem[63][0] ), .B(\u_div/PartRem[62][0] ), .Y(n7)
         );
  ADDHX1 U11 ( .A(\u_div/PartRem[2][4] ), .B(\u_div/u_add_PartRem_2_1/n3 ), 
        .CO(\u_div/u_add_PartRem_2_1/n2 ), .S(\u_div/SumTmp[1][4] ) );
  OR2X2 U12 ( .A(\u_div/PartRem[59][2] ), .B(\u_div/PartRem[59][3] ), .Y(
        \u_div/u_add_PartRem_2_58/n3 ) );
  NOR2BX4 U13 ( .AN(\u_div/PartRem[64][0] ), .B(n7), .Y(\u_div/CryTmp[59][6] )
         );
  XNOR2XL U14 ( .A(\u_div/PartRem[64][0] ), .B(n7), .Y(\u_div/SumTmp[59][4] )
         );
  XOR2XL U15 ( .A(\u_div/CryTmp[46][6] ), .B(n3), .Y(\u_div/QInv[46] ) );
  XOR2XL U16 ( .A(\u_div/CryTmp[47][6] ), .B(n4), .Y(\u_div/QInv[47] ) );
  XOR2XL U17 ( .A(\u_div/CryTmp[35][6] ), .B(n3), .Y(\u_div/QInv[35] ) );
  XOR2XL U18 ( .A(\u_div/CryTmp[36][6] ), .B(n4), .Y(\u_div/QInv[36] ) );
  XOR2XL U19 ( .A(\u_div/CryTmp[28][6] ), .B(n3), .Y(\u_div/QInv[28] ) );
  XOR2XL U20 ( .A(\u_div/CryTmp[25][6] ), .B(n3), .Y(\u_div/QInv[25] ) );
  XOR2XL U21 ( .A(\u_div/CryTmp[17][6] ), .B(n3), .Y(\u_div/QInv[17] ) );
  XOR2XL U22 ( .A(\u_div/CryTmp[6][6] ), .B(n4), .Y(\u_div/QInv[6] ) );
  XOR2XL U23 ( .A(\u_div/CryTmp[7][6] ), .B(n3), .Y(\u_div/QInv[7] ) );
  XOR2XL U24 ( .A(\u_div/CryTmp[53][6] ), .B(n2), .Y(\u_div/QInv[53] ) );
  XOR2XL U25 ( .A(\u_div/CryTmp[45][6] ), .B(n2), .Y(\u_div/QInv[45] ) );
  XOR2XL U26 ( .A(\u_div/CryTmp[48][6] ), .B(n2), .Y(\u_div/QInv[48] ) );
  INVXL U27 ( .A(\u_div/PartRem[59][2] ), .Y(\u_div/SumTmp[58][2] ) );
  INVXL U28 ( .A(\u_div/PartRem[3][2] ), .Y(\u_div/SumTmp[2][2] ) );
  INVX3 U29 ( .A(n1), .Y(n2) );
  ADDHX2 U30 ( .A(\u_div/PartRem[4][4] ), .B(\u_div/u_add_PartRem_2_3/n3 ), 
        .CO(\u_div/u_add_PartRem_2_3/n2 ), .S(\u_div/SumTmp[3][4] ) );
  OR2X2 U31 ( .A(\u_div/PartRem[4][2] ), .B(\u_div/PartRem[4][3] ), .Y(
        \u_div/u_add_PartRem_2_3/n3 ) );
  ADDHX2 U32 ( .A(\u_div/PartRem[59][4] ), .B(\u_div/u_add_PartRem_2_58/n3 ), 
        .CO(\u_div/u_add_PartRem_2_58/n2 ), .S(\u_div/SumTmp[58][4] ) );
  ADDHX2 U33 ( .A(\u_div/PartRem[53][4] ), .B(\u_div/u_add_PartRem_2_52/n3 ), 
        .CO(\u_div/u_add_PartRem_2_52/n2 ), .S(\u_div/SumTmp[52][4] ) );
  OR2X2 U34 ( .A(\u_div/PartRem[53][2] ), .B(\u_div/PartRem[53][3] ), .Y(
        \u_div/u_add_PartRem_2_52/n3 ) );
  ADDHX2 U35 ( .A(\u_div/PartRem[55][4] ), .B(\u_div/u_add_PartRem_2_54/n3 ), 
        .CO(\u_div/u_add_PartRem_2_54/n2 ), .S(\u_div/SumTmp[54][4] ) );
  OR2X2 U36 ( .A(\u_div/PartRem[55][2] ), .B(\u_div/PartRem[55][3] ), .Y(
        \u_div/u_add_PartRem_2_54/n3 ) );
  ADDHX2 U37 ( .A(\u_div/PartRem[48][4] ), .B(\u_div/u_add_PartRem_2_47/n3 ), 
        .CO(\u_div/u_add_PartRem_2_47/n2 ), .S(\u_div/SumTmp[47][4] ) );
  OR2X2 U38 ( .A(\u_div/PartRem[48][2] ), .B(\u_div/PartRem[48][3] ), .Y(
        \u_div/u_add_PartRem_2_47/n3 ) );
  ADDHX2 U39 ( .A(\u_div/PartRem[54][4] ), .B(\u_div/u_add_PartRem_2_53/n3 ), 
        .CO(\u_div/u_add_PartRem_2_53/n2 ), .S(\u_div/SumTmp[53][4] ) );
  OR2X2 U40 ( .A(\u_div/PartRem[54][2] ), .B(\u_div/PartRem[54][3] ), .Y(
        \u_div/u_add_PartRem_2_53/n3 ) );
  ADDHX2 U41 ( .A(\u_div/PartRem[45][4] ), .B(\u_div/u_add_PartRem_2_44/n3 ), 
        .CO(\u_div/u_add_PartRem_2_44/n2 ), .S(\u_div/SumTmp[44][4] ) );
  OR2X2 U42 ( .A(\u_div/PartRem[45][2] ), .B(\u_div/PartRem[45][3] ), .Y(
        \u_div/u_add_PartRem_2_44/n3 ) );
  OR2X2 U43 ( .A(\u_div/PartRem[52][2] ), .B(\u_div/PartRem[52][3] ), .Y(
        \u_div/u_add_PartRem_2_51/n3 ) );
  OR2X2 U44 ( .A(\u_div/PartRem[42][2] ), .B(\u_div/PartRem[42][3] ), .Y(
        \u_div/u_add_PartRem_2_41/n3 ) );
  OR2X2 U45 ( .A(\u_div/PartRem[47][2] ), .B(\u_div/PartRem[47][3] ), .Y(
        \u_div/u_add_PartRem_2_46/n3 ) );
  ADDHX2 U46 ( .A(\u_div/PartRem[44][4] ), .B(\u_div/u_add_PartRem_2_43/n3 ), 
        .CO(\u_div/u_add_PartRem_2_43/n2 ), .S(\u_div/SumTmp[43][4] ) );
  OR2X2 U47 ( .A(\u_div/PartRem[44][2] ), .B(\u_div/PartRem[44][3] ), .Y(
        \u_div/u_add_PartRem_2_43/n3 ) );
  ADDHX2 U48 ( .A(\u_div/PartRem[41][4] ), .B(\u_div/u_add_PartRem_2_40/n3 ), 
        .CO(\u_div/u_add_PartRem_2_40/n2 ), .S(\u_div/SumTmp[40][4] ) );
  OR2X2 U49 ( .A(\u_div/PartRem[41][2] ), .B(\u_div/PartRem[41][3] ), .Y(
        \u_div/u_add_PartRem_2_40/n3 ) );
  ADDHX2 U50 ( .A(\u_div/PartRem[51][4] ), .B(\u_div/u_add_PartRem_2_50/n3 ), 
        .CO(\u_div/u_add_PartRem_2_50/n2 ), .S(\u_div/SumTmp[50][4] ) );
  OR2X2 U51 ( .A(\u_div/PartRem[51][2] ), .B(\u_div/PartRem[51][3] ), .Y(
        \u_div/u_add_PartRem_2_50/n3 ) );
  ADDHX2 U52 ( .A(\u_div/PartRem[50][4] ), .B(\u_div/u_add_PartRem_2_49/n3 ), 
        .CO(\u_div/u_add_PartRem_2_49/n2 ), .S(\u_div/SumTmp[49][4] ) );
  OR2X2 U53 ( .A(\u_div/PartRem[50][2] ), .B(\u_div/PartRem[50][3] ), .Y(
        \u_div/u_add_PartRem_2_49/n3 ) );
  ADDHX2 U54 ( .A(\u_div/PartRem[49][4] ), .B(\u_div/u_add_PartRem_2_48/n3 ), 
        .CO(\u_div/u_add_PartRem_2_48/n2 ), .S(\u_div/SumTmp[48][4] ) );
  OR2X2 U55 ( .A(\u_div/PartRem[49][2] ), .B(\u_div/PartRem[49][3] ), .Y(
        \u_div/u_add_PartRem_2_48/n3 ) );
  ADDHX2 U56 ( .A(\u_div/PartRem[46][4] ), .B(\u_div/u_add_PartRem_2_45/n3 ), 
        .CO(\u_div/u_add_PartRem_2_45/n2 ), .S(\u_div/SumTmp[45][4] ) );
  OR2X2 U57 ( .A(\u_div/PartRem[46][2] ), .B(\u_div/PartRem[46][3] ), .Y(
        \u_div/u_add_PartRem_2_45/n3 ) );
  ADDHX2 U58 ( .A(\u_div/PartRem[43][4] ), .B(\u_div/u_add_PartRem_2_42/n3 ), 
        .CO(\u_div/u_add_PartRem_2_42/n2 ), .S(\u_div/SumTmp[42][4] ) );
  OR2X2 U59 ( .A(\u_div/PartRem[43][2] ), .B(\u_div/PartRem[43][3] ), .Y(
        \u_div/u_add_PartRem_2_42/n3 ) );
  ADDHX2 U60 ( .A(\u_div/PartRem[40][4] ), .B(\u_div/u_add_PartRem_2_39/n3 ), 
        .CO(\u_div/u_add_PartRem_2_39/n2 ), .S(\u_div/SumTmp[39][4] ) );
  OR2X2 U61 ( .A(\u_div/PartRem[40][2] ), .B(\u_div/PartRem[40][3] ), .Y(
        \u_div/u_add_PartRem_2_39/n3 ) );
  ADDHX2 U62 ( .A(\u_div/PartRem[39][4] ), .B(\u_div/u_add_PartRem_2_38/n3 ), 
        .CO(\u_div/u_add_PartRem_2_38/n2 ), .S(\u_div/SumTmp[38][4] ) );
  OR2X2 U63 ( .A(\u_div/PartRem[39][2] ), .B(\u_div/PartRem[39][3] ), .Y(
        \u_div/u_add_PartRem_2_38/n3 ) );
  OR2X2 U64 ( .A(\u_div/PartRem[37][2] ), .B(\u_div/PartRem[37][3] ), .Y(
        \u_div/u_add_PartRem_2_36/n3 ) );
  ADDHX2 U65 ( .A(\u_div/PartRem[36][4] ), .B(\u_div/u_add_PartRem_2_35/n3 ), 
        .CO(\u_div/u_add_PartRem_2_35/n2 ), .S(\u_div/SumTmp[35][4] ) );
  OR2X2 U66 ( .A(\u_div/PartRem[36][2] ), .B(\u_div/PartRem[36][3] ), .Y(
        \u_div/u_add_PartRem_2_35/n3 ) );
  ADDHX2 U67 ( .A(\u_div/PartRem[38][4] ), .B(\u_div/u_add_PartRem_2_37/n3 ), 
        .CO(\u_div/u_add_PartRem_2_37/n2 ), .S(\u_div/SumTmp[37][4] ) );
  OR2X2 U68 ( .A(\u_div/PartRem[38][2] ), .B(\u_div/PartRem[38][3] ), .Y(
        \u_div/u_add_PartRem_2_37/n3 ) );
  ADDHX2 U69 ( .A(\u_div/PartRem[35][4] ), .B(\u_div/u_add_PartRem_2_34/n3 ), 
        .CO(\u_div/u_add_PartRem_2_34/n2 ), .S(\u_div/SumTmp[34][4] ) );
  OR2X2 U70 ( .A(\u_div/PartRem[35][2] ), .B(\u_div/PartRem[35][3] ), .Y(
        \u_div/u_add_PartRem_2_34/n3 ) );
  ADDHX2 U71 ( .A(\u_div/PartRem[34][4] ), .B(\u_div/u_add_PartRem_2_33/n3 ), 
        .CO(\u_div/u_add_PartRem_2_33/n2 ), .S(\u_div/SumTmp[33][4] ) );
  OR2X2 U72 ( .A(\u_div/PartRem[34][2] ), .B(\u_div/PartRem[34][3] ), .Y(
        \u_div/u_add_PartRem_2_33/n3 ) );
  ADDHX2 U73 ( .A(\u_div/PartRem[15][4] ), .B(\u_div/u_add_PartRem_2_14/n3 ), 
        .CO(\u_div/u_add_PartRem_2_14/n2 ), .S(\u_div/SumTmp[14][4] ) );
  OR2X2 U74 ( .A(\u_div/PartRem[15][2] ), .B(\u_div/PartRem[15][3] ), .Y(
        \u_div/u_add_PartRem_2_14/n3 ) );
  ADDHX2 U75 ( .A(\u_div/PartRem[14][4] ), .B(\u_div/u_add_PartRem_2_13/n3 ), 
        .CO(\u_div/u_add_PartRem_2_13/n2 ), .S(\u_div/SumTmp[13][4] ) );
  OR2X2 U76 ( .A(\u_div/PartRem[14][2] ), .B(\u_div/PartRem[14][3] ), .Y(
        \u_div/u_add_PartRem_2_13/n3 ) );
  ADDHX2 U77 ( .A(\u_div/PartRem[16][4] ), .B(\u_div/u_add_PartRem_2_15/n3 ), 
        .CO(\u_div/u_add_PartRem_2_15/n2 ), .S(\u_div/SumTmp[15][4] ) );
  OR2X2 U78 ( .A(\u_div/PartRem[16][2] ), .B(\u_div/PartRem[16][3] ), .Y(
        \u_div/u_add_PartRem_2_15/n3 ) );
  ADDHX2 U79 ( .A(\u_div/PartRem[13][4] ), .B(\u_div/u_add_PartRem_2_12/n3 ), 
        .CO(\u_div/u_add_PartRem_2_12/n2 ), .S(\u_div/SumTmp[12][4] ) );
  OR2X2 U80 ( .A(\u_div/PartRem[13][2] ), .B(\u_div/PartRem[13][3] ), .Y(
        \u_div/u_add_PartRem_2_12/n3 ) );
  OR2X2 U81 ( .A(\u_div/PartRem[32][2] ), .B(\u_div/PartRem[32][3] ), .Y(
        \u_div/u_add_PartRem_2_31/n3 ) );
  ADDHX2 U82 ( .A(\u_div/PartRem[31][4] ), .B(\u_div/u_add_PartRem_2_30/n3 ), 
        .CO(\u_div/u_add_PartRem_2_30/n2 ), .S(\u_div/SumTmp[30][4] ) );
  OR2X2 U83 ( .A(\u_div/PartRem[31][2] ), .B(\u_div/PartRem[31][3] ), .Y(
        \u_div/u_add_PartRem_2_30/n3 ) );
  OR2X2 U84 ( .A(\u_div/PartRem[17][2] ), .B(\u_div/PartRem[17][3] ), .Y(
        \u_div/u_add_PartRem_2_16/n3 ) );
  ADDHX2 U85 ( .A(\u_div/PartRem[33][4] ), .B(\u_div/u_add_PartRem_2_32/n3 ), 
        .CO(\u_div/u_add_PartRem_2_32/n2 ), .S(\u_div/SumTmp[32][4] ) );
  OR2X2 U86 ( .A(\u_div/PartRem[33][2] ), .B(\u_div/PartRem[33][3] ), .Y(
        \u_div/u_add_PartRem_2_32/n3 ) );
  OR2X2 U87 ( .A(\u_div/PartRem[12][2] ), .B(\u_div/PartRem[12][3] ), .Y(
        \u_div/u_add_PartRem_2_11/n3 ) );
  ADDHX2 U88 ( .A(\u_div/PartRem[18][4] ), .B(\u_div/u_add_PartRem_2_17/n3 ), 
        .CO(\u_div/u_add_PartRem_2_17/n2 ), .S(\u_div/SumTmp[17][4] ) );
  OR2X2 U89 ( .A(\u_div/PartRem[18][2] ), .B(\u_div/PartRem[18][3] ), .Y(
        \u_div/u_add_PartRem_2_17/n3 ) );
  ADDHX2 U90 ( .A(\u_div/PartRem[30][4] ), .B(\u_div/u_add_PartRem_2_29/n3 ), 
        .CO(\u_div/u_add_PartRem_2_29/n2 ), .S(\u_div/SumTmp[29][4] ) );
  OR2X2 U91 ( .A(\u_div/PartRem[30][2] ), .B(\u_div/PartRem[30][3] ), .Y(
        \u_div/u_add_PartRem_2_29/n3 ) );
  ADDHX2 U92 ( .A(\u_div/PartRem[19][4] ), .B(\u_div/u_add_PartRem_2_18/n3 ), 
        .CO(\u_div/u_add_PartRem_2_18/n2 ), .S(\u_div/SumTmp[18][4] ) );
  OR2X2 U93 ( .A(\u_div/PartRem[19][2] ), .B(\u_div/PartRem[19][3] ), .Y(
        \u_div/u_add_PartRem_2_18/n3 ) );
  ADDHX2 U94 ( .A(\u_div/PartRem[29][4] ), .B(\u_div/u_add_PartRem_2_28/n3 ), 
        .CO(\u_div/u_add_PartRem_2_28/n2 ), .S(\u_div/SumTmp[28][4] ) );
  OR2X2 U95 ( .A(\u_div/PartRem[29][2] ), .B(\u_div/PartRem[29][3] ), .Y(
        \u_div/u_add_PartRem_2_28/n3 ) );
  ADDHX2 U96 ( .A(\u_div/PartRem[11][4] ), .B(\u_div/u_add_PartRem_2_10/n3 ), 
        .CO(\u_div/u_add_PartRem_2_10/n2 ), .S(\u_div/SumTmp[10][4] ) );
  OR2X2 U97 ( .A(\u_div/PartRem[11][2] ), .B(\u_div/PartRem[11][3] ), .Y(
        \u_div/u_add_PartRem_2_10/n3 ) );
  ADDHX2 U98 ( .A(\u_div/PartRem[20][4] ), .B(\u_div/u_add_PartRem_2_19/n3 ), 
        .CO(\u_div/u_add_PartRem_2_19/n2 ), .S(\u_div/SumTmp[19][4] ) );
  OR2X2 U99 ( .A(\u_div/PartRem[20][2] ), .B(\u_div/PartRem[20][3] ), .Y(
        \u_div/u_add_PartRem_2_19/n3 ) );
  ADDHX2 U100 ( .A(\u_div/PartRem[28][4] ), .B(\u_div/u_add_PartRem_2_27/n3 ), 
        .CO(\u_div/u_add_PartRem_2_27/n2 ), .S(\u_div/SumTmp[27][4] ) );
  OR2X2 U101 ( .A(\u_div/PartRem[28][2] ), .B(\u_div/PartRem[28][3] ), .Y(
        \u_div/u_add_PartRem_2_27/n3 ) );
  ADDHX2 U102 ( .A(\u_div/PartRem[21][4] ), .B(\u_div/u_add_PartRem_2_20/n3 ), 
        .CO(\u_div/u_add_PartRem_2_20/n2 ), .S(\u_div/SumTmp[20][4] ) );
  OR2X2 U103 ( .A(\u_div/PartRem[21][2] ), .B(\u_div/PartRem[21][3] ), .Y(
        \u_div/u_add_PartRem_2_20/n3 ) );
  ADDHX2 U104 ( .A(\u_div/PartRem[24][4] ), .B(\u_div/u_add_PartRem_2_23/n3 ), 
        .CO(\u_div/u_add_PartRem_2_23/n2 ), .S(\u_div/SumTmp[23][4] ) );
  OR2X2 U105 ( .A(\u_div/PartRem[24][2] ), .B(\u_div/PartRem[24][3] ), .Y(
        \u_div/u_add_PartRem_2_23/n3 ) );
  ADDHX2 U106 ( .A(\u_div/PartRem[26][4] ), .B(\u_div/u_add_PartRem_2_25/n3 ), 
        .CO(\u_div/u_add_PartRem_2_25/n2 ), .S(\u_div/SumTmp[25][4] ) );
  OR2X2 U107 ( .A(\u_div/PartRem[26][2] ), .B(\u_div/PartRem[26][3] ), .Y(
        \u_div/u_add_PartRem_2_25/n3 ) );
  ADDHX2 U108 ( .A(\u_div/PartRem[23][4] ), .B(\u_div/u_add_PartRem_2_22/n3 ), 
        .CO(\u_div/u_add_PartRem_2_22/n2 ), .S(\u_div/SumTmp[22][4] ) );
  OR2X2 U109 ( .A(\u_div/PartRem[23][2] ), .B(\u_div/PartRem[23][3] ), .Y(
        \u_div/u_add_PartRem_2_22/n3 ) );
  ADDHX2 U110 ( .A(\u_div/PartRem[25][4] ), .B(\u_div/u_add_PartRem_2_24/n3 ), 
        .CO(\u_div/u_add_PartRem_2_24/n2 ), .S(\u_div/SumTmp[24][4] ) );
  OR2X2 U111 ( .A(\u_div/PartRem[25][2] ), .B(\u_div/PartRem[25][3] ), .Y(
        \u_div/u_add_PartRem_2_24/n3 ) );
  ADDHX2 U112 ( .A(\u_div/PartRem[8][4] ), .B(\u_div/u_add_PartRem_2_7/n3 ), 
        .CO(\u_div/u_add_PartRem_2_7/n2 ), .S(\u_div/SumTmp[7][4] ) );
  OR2X2 U113 ( .A(\u_div/PartRem[8][2] ), .B(\u_div/PartRem[8][3] ), .Y(
        \u_div/u_add_PartRem_2_7/n3 ) );
  ADDHX2 U114 ( .A(\u_div/PartRem[9][4] ), .B(\u_div/u_add_PartRem_2_8/n3 ), 
        .CO(\u_div/u_add_PartRem_2_8/n2 ), .S(\u_div/SumTmp[8][4] ) );
  OR2X2 U115 ( .A(\u_div/PartRem[9][2] ), .B(\u_div/PartRem[9][3] ), .Y(
        \u_div/u_add_PartRem_2_8/n3 ) );
  ADDHX2 U116 ( .A(\u_div/PartRem[10][4] ), .B(\u_div/u_add_PartRem_2_9/n3 ), 
        .CO(\u_div/u_add_PartRem_2_9/n2 ), .S(\u_div/SumTmp[9][4] ) );
  OR2X2 U117 ( .A(\u_div/PartRem[10][2] ), .B(\u_div/PartRem[10][3] ), .Y(
        \u_div/u_add_PartRem_2_9/n3 ) );
  ADDHX2 U118 ( .A(\u_div/PartRem[6][4] ), .B(\u_div/u_add_PartRem_2_5/n3 ), 
        .CO(\u_div/u_add_PartRem_2_5/n2 ), .S(\u_div/SumTmp[5][4] ) );
  OR2X2 U119 ( .A(\u_div/PartRem[6][2] ), .B(\u_div/PartRem[6][3] ), .Y(
        \u_div/u_add_PartRem_2_5/n3 ) );
  ADDHX2 U120 ( .A(\u_div/PartRem[5][4] ), .B(\u_div/u_add_PartRem_2_4/n3 ), 
        .CO(\u_div/u_add_PartRem_2_4/n2 ), .S(\u_div/SumTmp[4][4] ) );
  OR2X2 U121 ( .A(\u_div/PartRem[5][2] ), .B(\u_div/PartRem[5][3] ), .Y(
        \u_div/u_add_PartRem_2_4/n3 ) );
  OR2X2 U122 ( .A(\u_div/PartRem[2][2] ), .B(\u_div/PartRem[2][3] ), .Y(
        \u_div/u_add_PartRem_2_1/n3 ) );
  ADDHX2 U123 ( .A(\u_div/PartRem[58][4] ), .B(\u_div/u_add_PartRem_2_57/n3 ), 
        .CO(\u_div/u_add_PartRem_2_57/n2 ), .S(\u_div/SumTmp[57][4] ) );
  OR2X2 U124 ( .A(\u_div/PartRem[58][2] ), .B(\u_div/PartRem[58][3] ), .Y(
        \u_div/u_add_PartRem_2_57/n3 ) );
  ADDHX2 U125 ( .A(\u_div/PartRem[56][4] ), .B(\u_div/u_add_PartRem_2_55/n3 ), 
        .CO(\u_div/u_add_PartRem_2_55/n2 ), .S(\u_div/SumTmp[55][4] ) );
  OR2X2 U126 ( .A(\u_div/PartRem[56][2] ), .B(\u_div/PartRem[56][3] ), .Y(
        \u_div/u_add_PartRem_2_55/n3 ) );
  OR2X2 U127 ( .A(\u_div/PartRem[57][2] ), .B(\u_div/PartRem[57][3] ), .Y(
        \u_div/u_add_PartRem_2_56/n3 ) );
  OR2X4 U128 ( .A(\u_div/PartRem[1][3] ), .B(\u_div/PartRem[1][2] ), .Y(n5) );
  INVXL U129 ( .A(\u_div/PartRem[2][2] ), .Y(\u_div/SumTmp[1][2] ) );
  OR2X1 U130 ( .A(\u_div/PartRem[2][5] ), .B(\u_div/u_add_PartRem_2_1/n2 ), 
        .Y(\u_div/CryTmp[1][6] ) );
  XOR2X1 U131 ( .A(\u_div/CryTmp[0][6] ), .B(n4), .Y(\u_div/QInv[0] ) );
  AO21X1 U132 ( .A0(\u_div/PartRem[1][4] ), .A1(n5), .B0(\u_div/PartRem[1][5] ), .Y(\u_div/CryTmp[0][6] ) );
  MXI2X1 U133 ( .A(n6), .B(\u_div/PartRem[62][0] ), .S0(\u_div/CryTmp[59][6] ), 
        .Y(\u_div/PartRem[59][3] ) );
  CLKINVX1 U134 ( .A(\u_div/PartRem[62][0] ), .Y(n6) );
  MXI2X1 U135 ( .A(\u_div/SumTmp[22][2] ), .B(\u_div/PartRem[23][2] ), .S0(
        \u_div/CryTmp[22][6] ), .Y(\u_div/PartRem[22][3] ) );
  CLKINVX1 U136 ( .A(\u_div/PartRem[23][2] ), .Y(\u_div/SumTmp[22][2] ) );
  MXI2X1 U137 ( .A(\u_div/SumTmp[12][2] ), .B(\u_div/PartRem[13][2] ), .S0(
        \u_div/CryTmp[12][6] ), .Y(\u_div/PartRem[12][3] ) );
  CLKINVX1 U138 ( .A(\u_div/PartRem[13][2] ), .Y(\u_div/SumTmp[12][2] ) );
  MXI2X1 U139 ( .A(\u_div/SumTmp[57][2] ), .B(\u_div/PartRem[58][2] ), .S0(
        \u_div/CryTmp[57][6] ), .Y(\u_div/PartRem[57][3] ) );
  CLKINVX1 U140 ( .A(\u_div/PartRem[58][2] ), .Y(\u_div/SumTmp[57][2] ) );
  MXI2X1 U141 ( .A(\u_div/SumTmp[52][2] ), .B(\u_div/PartRem[53][2] ), .S0(
        \u_div/CryTmp[52][6] ), .Y(\u_div/PartRem[52][3] ) );
  CLKINVX1 U142 ( .A(\u_div/PartRem[53][2] ), .Y(\u_div/SumTmp[52][2] ) );
  MXI2X1 U143 ( .A(\u_div/SumTmp[47][2] ), .B(\u_div/PartRem[48][2] ), .S0(
        \u_div/CryTmp[47][6] ), .Y(\u_div/PartRem[47][3] ) );
  CLKINVX1 U144 ( .A(\u_div/PartRem[48][2] ), .Y(\u_div/SumTmp[47][2] ) );
  MXI2X1 U145 ( .A(\u_div/SumTmp[42][2] ), .B(\u_div/PartRem[43][2] ), .S0(
        \u_div/CryTmp[42][6] ), .Y(\u_div/PartRem[42][3] ) );
  CLKINVX1 U146 ( .A(\u_div/PartRem[43][2] ), .Y(\u_div/SumTmp[42][2] ) );
  MXI2X1 U147 ( .A(\u_div/SumTmp[37][2] ), .B(\u_div/PartRem[38][2] ), .S0(
        \u_div/CryTmp[37][6] ), .Y(\u_div/PartRem[37][3] ) );
  CLKINVX1 U148 ( .A(\u_div/PartRem[38][2] ), .Y(\u_div/SumTmp[37][2] ) );
  MXI2X1 U149 ( .A(\u_div/SumTmp[32][2] ), .B(\u_div/PartRem[33][2] ), .S0(
        \u_div/CryTmp[32][6] ), .Y(\u_div/PartRem[32][3] ) );
  CLKINVX1 U150 ( .A(\u_div/PartRem[33][2] ), .Y(\u_div/SumTmp[32][2] ) );
  MXI2X1 U151 ( .A(\u_div/SumTmp[27][2] ), .B(\u_div/PartRem[28][2] ), .S0(
        \u_div/CryTmp[27][6] ), .Y(\u_div/PartRem[27][3] ) );
  CLKINVX1 U152 ( .A(\u_div/PartRem[28][2] ), .Y(\u_div/SumTmp[27][2] ) );
  MXI2X1 U153 ( .A(\u_div/SumTmp[17][2] ), .B(\u_div/PartRem[18][2] ), .S0(
        \u_div/CryTmp[17][6] ), .Y(\u_div/PartRem[17][3] ) );
  CLKINVX1 U154 ( .A(\u_div/PartRem[18][2] ), .Y(\u_div/SumTmp[17][2] ) );
  MXI2X1 U155 ( .A(\u_div/SumTmp[7][2] ), .B(\u_div/PartRem[8][2] ), .S0(
        \u_div/CryTmp[7][6] ), .Y(\u_div/PartRem[7][3] ) );
  CLKINVX1 U156 ( .A(\u_div/PartRem[8][2] ), .Y(\u_div/SumTmp[7][2] ) );
  MXI2X1 U157 ( .A(\u_div/SumTmp[58][2] ), .B(\u_div/PartRem[59][2] ), .S0(
        \u_div/CryTmp[58][6] ), .Y(\u_div/PartRem[58][3] ) );
  MXI2X1 U158 ( .A(\u_div/SumTmp[56][2] ), .B(\u_div/PartRem[57][2] ), .S0(
        \u_div/CryTmp[56][6] ), .Y(\u_div/PartRem[56][3] ) );
  CLKINVX1 U159 ( .A(\u_div/PartRem[57][2] ), .Y(\u_div/SumTmp[56][2] ) );
  MXI2X1 U160 ( .A(\u_div/SumTmp[55][2] ), .B(\u_div/PartRem[56][2] ), .S0(
        \u_div/CryTmp[55][6] ), .Y(\u_div/PartRem[55][3] ) );
  CLKINVX1 U161 ( .A(\u_div/PartRem[56][2] ), .Y(\u_div/SumTmp[55][2] ) );
  MXI2X1 U162 ( .A(\u_div/SumTmp[54][2] ), .B(\u_div/PartRem[55][2] ), .S0(
        \u_div/CryTmp[54][6] ), .Y(\u_div/PartRem[54][3] ) );
  CLKINVX1 U163 ( .A(\u_div/PartRem[55][2] ), .Y(\u_div/SumTmp[54][2] ) );
  MXI2X1 U164 ( .A(\u_div/SumTmp[53][2] ), .B(\u_div/PartRem[54][2] ), .S0(
        \u_div/CryTmp[53][6] ), .Y(\u_div/PartRem[53][3] ) );
  CLKINVX1 U165 ( .A(\u_div/PartRem[54][2] ), .Y(\u_div/SumTmp[53][2] ) );
  MXI2X1 U166 ( .A(\u_div/SumTmp[51][2] ), .B(\u_div/PartRem[52][2] ), .S0(
        \u_div/CryTmp[51][6] ), .Y(\u_div/PartRem[51][3] ) );
  CLKINVX1 U167 ( .A(\u_div/PartRem[52][2] ), .Y(\u_div/SumTmp[51][2] ) );
  MXI2X1 U168 ( .A(\u_div/SumTmp[50][2] ), .B(\u_div/PartRem[51][2] ), .S0(
        \u_div/CryTmp[50][6] ), .Y(\u_div/PartRem[50][3] ) );
  CLKINVX1 U169 ( .A(\u_div/PartRem[51][2] ), .Y(\u_div/SumTmp[50][2] ) );
  MXI2X1 U170 ( .A(\u_div/SumTmp[49][2] ), .B(\u_div/PartRem[50][2] ), .S0(
        \u_div/CryTmp[49][6] ), .Y(\u_div/PartRem[49][3] ) );
  CLKINVX1 U171 ( .A(\u_div/PartRem[50][2] ), .Y(\u_div/SumTmp[49][2] ) );
  MXI2X1 U172 ( .A(\u_div/SumTmp[48][2] ), .B(\u_div/PartRem[49][2] ), .S0(
        \u_div/CryTmp[48][6] ), .Y(\u_div/PartRem[48][3] ) );
  CLKINVX1 U173 ( .A(\u_div/PartRem[49][2] ), .Y(\u_div/SumTmp[48][2] ) );
  MXI2X1 U174 ( .A(\u_div/SumTmp[46][2] ), .B(\u_div/PartRem[47][2] ), .S0(
        \u_div/CryTmp[46][6] ), .Y(\u_div/PartRem[46][3] ) );
  CLKINVX1 U175 ( .A(\u_div/PartRem[47][2] ), .Y(\u_div/SumTmp[46][2] ) );
  MXI2X1 U176 ( .A(\u_div/SumTmp[45][2] ), .B(\u_div/PartRem[46][2] ), .S0(
        \u_div/CryTmp[45][6] ), .Y(\u_div/PartRem[45][3] ) );
  CLKINVX1 U177 ( .A(\u_div/PartRem[46][2] ), .Y(\u_div/SumTmp[45][2] ) );
  MXI2X1 U178 ( .A(\u_div/SumTmp[44][2] ), .B(\u_div/PartRem[45][2] ), .S0(
        \u_div/CryTmp[44][6] ), .Y(\u_div/PartRem[44][3] ) );
  CLKINVX1 U179 ( .A(\u_div/PartRem[45][2] ), .Y(\u_div/SumTmp[44][2] ) );
  MXI2X1 U180 ( .A(\u_div/SumTmp[43][2] ), .B(\u_div/PartRem[44][2] ), .S0(
        \u_div/CryTmp[43][6] ), .Y(\u_div/PartRem[43][3] ) );
  CLKINVX1 U181 ( .A(\u_div/PartRem[44][2] ), .Y(\u_div/SumTmp[43][2] ) );
  MXI2X1 U182 ( .A(\u_div/SumTmp[41][2] ), .B(\u_div/PartRem[42][2] ), .S0(
        \u_div/CryTmp[41][6] ), .Y(\u_div/PartRem[41][3] ) );
  CLKINVX1 U183 ( .A(\u_div/PartRem[42][2] ), .Y(\u_div/SumTmp[41][2] ) );
  MXI2X1 U184 ( .A(\u_div/SumTmp[40][2] ), .B(\u_div/PartRem[41][2] ), .S0(
        \u_div/CryTmp[40][6] ), .Y(\u_div/PartRem[40][3] ) );
  CLKINVX1 U185 ( .A(\u_div/PartRem[41][2] ), .Y(\u_div/SumTmp[40][2] ) );
  MXI2X1 U186 ( .A(\u_div/SumTmp[39][2] ), .B(\u_div/PartRem[40][2] ), .S0(
        \u_div/CryTmp[39][6] ), .Y(\u_div/PartRem[39][3] ) );
  CLKINVX1 U187 ( .A(\u_div/PartRem[40][2] ), .Y(\u_div/SumTmp[39][2] ) );
  MXI2X1 U188 ( .A(\u_div/SumTmp[38][2] ), .B(\u_div/PartRem[39][2] ), .S0(
        \u_div/CryTmp[38][6] ), .Y(\u_div/PartRem[38][3] ) );
  CLKINVX1 U189 ( .A(\u_div/PartRem[39][2] ), .Y(\u_div/SumTmp[38][2] ) );
  MXI2X1 U190 ( .A(\u_div/SumTmp[36][2] ), .B(\u_div/PartRem[37][2] ), .S0(
        \u_div/CryTmp[36][6] ), .Y(\u_div/PartRem[36][3] ) );
  CLKINVX1 U191 ( .A(\u_div/PartRem[37][2] ), .Y(\u_div/SumTmp[36][2] ) );
  MXI2X1 U192 ( .A(\u_div/SumTmp[35][2] ), .B(\u_div/PartRem[36][2] ), .S0(
        \u_div/CryTmp[35][6] ), .Y(\u_div/PartRem[35][3] ) );
  CLKINVX1 U193 ( .A(\u_div/PartRem[36][2] ), .Y(\u_div/SumTmp[35][2] ) );
  MXI2X1 U194 ( .A(\u_div/SumTmp[34][2] ), .B(\u_div/PartRem[35][2] ), .S0(
        \u_div/CryTmp[34][6] ), .Y(\u_div/PartRem[34][3] ) );
  CLKINVX1 U195 ( .A(\u_div/PartRem[35][2] ), .Y(\u_div/SumTmp[34][2] ) );
  MXI2X1 U196 ( .A(\u_div/SumTmp[33][2] ), .B(\u_div/PartRem[34][2] ), .S0(
        \u_div/CryTmp[33][6] ), .Y(\u_div/PartRem[33][3] ) );
  CLKINVX1 U197 ( .A(\u_div/PartRem[34][2] ), .Y(\u_div/SumTmp[33][2] ) );
  MXI2X1 U198 ( .A(\u_div/SumTmp[31][2] ), .B(\u_div/PartRem[32][2] ), .S0(
        \u_div/CryTmp[31][6] ), .Y(\u_div/PartRem[31][3] ) );
  CLKINVX1 U199 ( .A(\u_div/PartRem[32][2] ), .Y(\u_div/SumTmp[31][2] ) );
  MXI2X1 U200 ( .A(\u_div/SumTmp[30][2] ), .B(\u_div/PartRem[31][2] ), .S0(
        \u_div/CryTmp[30][6] ), .Y(\u_div/PartRem[30][3] ) );
  CLKINVX1 U201 ( .A(\u_div/PartRem[31][2] ), .Y(\u_div/SumTmp[30][2] ) );
  MXI2X1 U202 ( .A(\u_div/SumTmp[29][2] ), .B(\u_div/PartRem[30][2] ), .S0(
        \u_div/CryTmp[29][6] ), .Y(\u_div/PartRem[29][3] ) );
  CLKINVX1 U203 ( .A(\u_div/PartRem[30][2] ), .Y(\u_div/SumTmp[29][2] ) );
  MXI2X1 U204 ( .A(\u_div/SumTmp[28][2] ), .B(\u_div/PartRem[29][2] ), .S0(
        \u_div/CryTmp[28][6] ), .Y(\u_div/PartRem[28][3] ) );
  CLKINVX1 U205 ( .A(\u_div/PartRem[29][2] ), .Y(\u_div/SumTmp[28][2] ) );
  MXI2X1 U206 ( .A(\u_div/SumTmp[26][2] ), .B(\u_div/PartRem[27][2] ), .S0(
        \u_div/CryTmp[26][6] ), .Y(\u_div/PartRem[26][3] ) );
  CLKINVX1 U207 ( .A(\u_div/PartRem[27][2] ), .Y(\u_div/SumTmp[26][2] ) );
  MXI2X1 U208 ( .A(\u_div/SumTmp[25][2] ), .B(\u_div/PartRem[26][2] ), .S0(
        \u_div/CryTmp[25][6] ), .Y(\u_div/PartRem[25][3] ) );
  CLKINVX1 U209 ( .A(\u_div/PartRem[26][2] ), .Y(\u_div/SumTmp[25][2] ) );
  MXI2X1 U210 ( .A(\u_div/SumTmp[24][2] ), .B(\u_div/PartRem[25][2] ), .S0(
        \u_div/CryTmp[24][6] ), .Y(\u_div/PartRem[24][3] ) );
  CLKINVX1 U211 ( .A(\u_div/PartRem[25][2] ), .Y(\u_div/SumTmp[24][2] ) );
  MXI2X1 U212 ( .A(\u_div/SumTmp[23][2] ), .B(\u_div/PartRem[24][2] ), .S0(
        \u_div/CryTmp[23][6] ), .Y(\u_div/PartRem[23][3] ) );
  CLKINVX1 U213 ( .A(\u_div/PartRem[24][2] ), .Y(\u_div/SumTmp[23][2] ) );
  MXI2X1 U214 ( .A(\u_div/SumTmp[21][2] ), .B(\u_div/PartRem[22][2] ), .S0(
        \u_div/CryTmp[21][6] ), .Y(\u_div/PartRem[21][3] ) );
  CLKINVX1 U215 ( .A(\u_div/PartRem[22][2] ), .Y(\u_div/SumTmp[21][2] ) );
  MXI2X1 U216 ( .A(\u_div/SumTmp[20][2] ), .B(\u_div/PartRem[21][2] ), .S0(
        \u_div/CryTmp[20][6] ), .Y(\u_div/PartRem[20][3] ) );
  CLKINVX1 U217 ( .A(\u_div/PartRem[21][2] ), .Y(\u_div/SumTmp[20][2] ) );
  MXI2X1 U218 ( .A(\u_div/SumTmp[19][2] ), .B(\u_div/PartRem[20][2] ), .S0(
        \u_div/CryTmp[19][6] ), .Y(\u_div/PartRem[19][3] ) );
  CLKINVX1 U219 ( .A(\u_div/PartRem[20][2] ), .Y(\u_div/SumTmp[19][2] ) );
  MXI2X1 U220 ( .A(\u_div/SumTmp[18][2] ), .B(\u_div/PartRem[19][2] ), .S0(
        \u_div/CryTmp[18][6] ), .Y(\u_div/PartRem[18][3] ) );
  CLKINVX1 U221 ( .A(\u_div/PartRem[19][2] ), .Y(\u_div/SumTmp[18][2] ) );
  MXI2X1 U222 ( .A(\u_div/SumTmp[16][2] ), .B(\u_div/PartRem[17][2] ), .S0(
        \u_div/CryTmp[16][6] ), .Y(\u_div/PartRem[16][3] ) );
  CLKINVX1 U223 ( .A(\u_div/PartRem[17][2] ), .Y(\u_div/SumTmp[16][2] ) );
  MXI2X1 U224 ( .A(\u_div/SumTmp[15][2] ), .B(\u_div/PartRem[16][2] ), .S0(
        \u_div/CryTmp[15][6] ), .Y(\u_div/PartRem[15][3] ) );
  CLKINVX1 U225 ( .A(\u_div/PartRem[16][2] ), .Y(\u_div/SumTmp[15][2] ) );
  MXI2X1 U226 ( .A(\u_div/SumTmp[14][2] ), .B(\u_div/PartRem[15][2] ), .S0(
        \u_div/CryTmp[14][6] ), .Y(\u_div/PartRem[14][3] ) );
  CLKINVX1 U227 ( .A(\u_div/PartRem[15][2] ), .Y(\u_div/SumTmp[14][2] ) );
  MXI2X1 U228 ( .A(\u_div/SumTmp[13][2] ), .B(\u_div/PartRem[14][2] ), .S0(
        \u_div/CryTmp[13][6] ), .Y(\u_div/PartRem[13][3] ) );
  CLKINVX1 U229 ( .A(\u_div/PartRem[14][2] ), .Y(\u_div/SumTmp[13][2] ) );
  MXI2X1 U230 ( .A(\u_div/SumTmp[11][2] ), .B(\u_div/PartRem[12][2] ), .S0(
        \u_div/CryTmp[11][6] ), .Y(\u_div/PartRem[11][3] ) );
  CLKINVX1 U231 ( .A(\u_div/PartRem[12][2] ), .Y(\u_div/SumTmp[11][2] ) );
  MXI2X1 U232 ( .A(\u_div/SumTmp[10][2] ), .B(\u_div/PartRem[11][2] ), .S0(
        \u_div/CryTmp[10][6] ), .Y(\u_div/PartRem[10][3] ) );
  CLKINVX1 U233 ( .A(\u_div/PartRem[11][2] ), .Y(\u_div/SumTmp[10][2] ) );
  MXI2X1 U234 ( .A(\u_div/SumTmp[9][2] ), .B(\u_div/PartRem[10][2] ), .S0(
        \u_div/CryTmp[9][6] ), .Y(\u_div/PartRem[9][3] ) );
  CLKINVX1 U235 ( .A(\u_div/PartRem[10][2] ), .Y(\u_div/SumTmp[9][2] ) );
  MXI2X1 U236 ( .A(\u_div/SumTmp[8][2] ), .B(\u_div/PartRem[9][2] ), .S0(
        \u_div/CryTmp[8][6] ), .Y(\u_div/PartRem[8][3] ) );
  CLKINVX1 U237 ( .A(\u_div/PartRem[9][2] ), .Y(\u_div/SumTmp[8][2] ) );
  MXI2X1 U238 ( .A(\u_div/SumTmp[6][2] ), .B(\u_div/PartRem[7][2] ), .S0(
        \u_div/CryTmp[6][6] ), .Y(\u_div/PartRem[6][3] ) );
  CLKINVX1 U239 ( .A(\u_div/PartRem[7][2] ), .Y(\u_div/SumTmp[6][2] ) );
  MXI2X1 U240 ( .A(\u_div/SumTmp[5][2] ), .B(\u_div/PartRem[6][2] ), .S0(
        \u_div/CryTmp[5][6] ), .Y(\u_div/PartRem[5][3] ) );
  CLKINVX1 U241 ( .A(\u_div/PartRem[6][2] ), .Y(\u_div/SumTmp[5][2] ) );
  MXI2X1 U242 ( .A(\u_div/SumTmp[4][2] ), .B(\u_div/PartRem[5][2] ), .S0(
        \u_div/CryTmp[4][6] ), .Y(\u_div/PartRem[4][3] ) );
  CLKINVX1 U243 ( .A(\u_div/PartRem[5][2] ), .Y(\u_div/SumTmp[4][2] ) );
  MXI2X1 U244 ( .A(\u_div/SumTmp[2][2] ), .B(\u_div/PartRem[3][2] ), .S0(
        \u_div/CryTmp[2][6] ), .Y(\u_div/PartRem[2][3] ) );
  CLKINVX1 U245 ( .A(\u_div/PartRem[4][2] ), .Y(\u_div/SumTmp[3][2] ) );
  INVX4 U246 ( .A(n1), .Y(n4) );
  INVX4 U247 ( .A(n1), .Y(n3) );
  OR2X2 U248 ( .A(\u_div/PartRem[4][5] ), .B(\u_div/u_add_PartRem_2_3/n2 ), 
        .Y(\u_div/CryTmp[3][6] ) );
  OR2X1 U249 ( .A(\u_div/PartRem[59][5] ), .B(\u_div/u_add_PartRem_2_58/n2 ), 
        .Y(\u_div/CryTmp[58][6] ) );
  XNOR2X1 U250 ( .A(\u_div/PartRem[59][3] ), .B(\u_div/PartRem[59][2] ), .Y(
        \u_div/SumTmp[58][3] ) );
  OR2X1 U251 ( .A(\u_div/PartRem[58][5] ), .B(\u_div/u_add_PartRem_2_57/n2 ), 
        .Y(\u_div/CryTmp[57][6] ) );
  XNOR2X1 U252 ( .A(\u_div/PartRem[58][3] ), .B(\u_div/PartRem[58][2] ), .Y(
        \u_div/SumTmp[57][3] ) );
  OR2X1 U253 ( .A(\u_div/PartRem[57][5] ), .B(\u_div/u_add_PartRem_2_56/n2 ), 
        .Y(\u_div/CryTmp[56][6] ) );
  XNOR2X1 U254 ( .A(\u_div/PartRem[57][3] ), .B(\u_div/PartRem[57][2] ), .Y(
        \u_div/SumTmp[56][3] ) );
  OR2X1 U255 ( .A(\u_div/PartRem[56][5] ), .B(\u_div/u_add_PartRem_2_55/n2 ), 
        .Y(\u_div/CryTmp[55][6] ) );
  XNOR2X1 U256 ( .A(\u_div/PartRem[56][3] ), .B(\u_div/PartRem[56][2] ), .Y(
        \u_div/SumTmp[55][3] ) );
  OR2X1 U257 ( .A(\u_div/PartRem[55][5] ), .B(\u_div/u_add_PartRem_2_54/n2 ), 
        .Y(\u_div/CryTmp[54][6] ) );
  XNOR2X1 U258 ( .A(\u_div/PartRem[55][3] ), .B(\u_div/PartRem[55][2] ), .Y(
        \u_div/SumTmp[54][3] ) );
  OR2X1 U259 ( .A(\u_div/PartRem[54][5] ), .B(\u_div/u_add_PartRem_2_53/n2 ), 
        .Y(\u_div/CryTmp[53][6] ) );
  XNOR2X1 U260 ( .A(\u_div/PartRem[54][3] ), .B(\u_div/PartRem[54][2] ), .Y(
        \u_div/SumTmp[53][3] ) );
  OR2X1 U261 ( .A(\u_div/PartRem[53][5] ), .B(\u_div/u_add_PartRem_2_52/n2 ), 
        .Y(\u_div/CryTmp[52][6] ) );
  XNOR2X1 U262 ( .A(\u_div/PartRem[53][3] ), .B(\u_div/PartRem[53][2] ), .Y(
        \u_div/SumTmp[52][3] ) );
  OR2X1 U263 ( .A(\u_div/PartRem[52][5] ), .B(\u_div/u_add_PartRem_2_51/n2 ), 
        .Y(\u_div/CryTmp[51][6] ) );
  XNOR2X1 U264 ( .A(\u_div/PartRem[52][3] ), .B(\u_div/PartRem[52][2] ), .Y(
        \u_div/SumTmp[51][3] ) );
  OR2X1 U265 ( .A(\u_div/PartRem[51][5] ), .B(\u_div/u_add_PartRem_2_50/n2 ), 
        .Y(\u_div/CryTmp[50][6] ) );
  XNOR2X1 U266 ( .A(\u_div/PartRem[51][3] ), .B(\u_div/PartRem[51][2] ), .Y(
        \u_div/SumTmp[50][3] ) );
  OR2X1 U267 ( .A(\u_div/PartRem[50][5] ), .B(\u_div/u_add_PartRem_2_49/n2 ), 
        .Y(\u_div/CryTmp[49][6] ) );
  XNOR2X1 U268 ( .A(\u_div/PartRem[50][3] ), .B(\u_div/PartRem[50][2] ), .Y(
        \u_div/SumTmp[49][3] ) );
  OR2X1 U269 ( .A(\u_div/PartRem[49][5] ), .B(\u_div/u_add_PartRem_2_48/n2 ), 
        .Y(\u_div/CryTmp[48][6] ) );
  XNOR2X1 U270 ( .A(\u_div/PartRem[49][3] ), .B(\u_div/PartRem[49][2] ), .Y(
        \u_div/SumTmp[48][3] ) );
  OR2X1 U271 ( .A(\u_div/PartRem[48][5] ), .B(\u_div/u_add_PartRem_2_47/n2 ), 
        .Y(\u_div/CryTmp[47][6] ) );
  XNOR2X1 U272 ( .A(\u_div/PartRem[48][3] ), .B(\u_div/PartRem[48][2] ), .Y(
        \u_div/SumTmp[47][3] ) );
  OR2X1 U273 ( .A(\u_div/PartRem[47][5] ), .B(\u_div/u_add_PartRem_2_46/n2 ), 
        .Y(\u_div/CryTmp[46][6] ) );
  XNOR2X1 U274 ( .A(\u_div/PartRem[47][3] ), .B(\u_div/PartRem[47][2] ), .Y(
        \u_div/SumTmp[46][3] ) );
  OR2X1 U275 ( .A(\u_div/PartRem[46][5] ), .B(\u_div/u_add_PartRem_2_45/n2 ), 
        .Y(\u_div/CryTmp[45][6] ) );
  XNOR2X1 U276 ( .A(\u_div/PartRem[46][3] ), .B(\u_div/PartRem[46][2] ), .Y(
        \u_div/SumTmp[45][3] ) );
  OR2X1 U277 ( .A(\u_div/PartRem[45][5] ), .B(\u_div/u_add_PartRem_2_44/n2 ), 
        .Y(\u_div/CryTmp[44][6] ) );
  XNOR2X1 U278 ( .A(\u_div/PartRem[45][3] ), .B(\u_div/PartRem[45][2] ), .Y(
        \u_div/SumTmp[44][3] ) );
  OR2X1 U279 ( .A(\u_div/PartRem[44][5] ), .B(\u_div/u_add_PartRem_2_43/n2 ), 
        .Y(\u_div/CryTmp[43][6] ) );
  XNOR2X1 U280 ( .A(\u_div/PartRem[44][3] ), .B(\u_div/PartRem[44][2] ), .Y(
        \u_div/SumTmp[43][3] ) );
  OR2X1 U281 ( .A(\u_div/PartRem[43][5] ), .B(\u_div/u_add_PartRem_2_42/n2 ), 
        .Y(\u_div/CryTmp[42][6] ) );
  XNOR2X1 U282 ( .A(\u_div/PartRem[43][3] ), .B(\u_div/PartRem[43][2] ), .Y(
        \u_div/SumTmp[42][3] ) );
  OR2X1 U283 ( .A(\u_div/PartRem[42][5] ), .B(\u_div/u_add_PartRem_2_41/n2 ), 
        .Y(\u_div/CryTmp[41][6] ) );
  XNOR2X1 U284 ( .A(\u_div/PartRem[42][3] ), .B(\u_div/PartRem[42][2] ), .Y(
        \u_div/SumTmp[41][3] ) );
  OR2X1 U285 ( .A(\u_div/PartRem[41][5] ), .B(\u_div/u_add_PartRem_2_40/n2 ), 
        .Y(\u_div/CryTmp[40][6] ) );
  XNOR2X1 U286 ( .A(\u_div/PartRem[41][3] ), .B(\u_div/PartRem[41][2] ), .Y(
        \u_div/SumTmp[40][3] ) );
  OR2X1 U287 ( .A(\u_div/PartRem[40][5] ), .B(\u_div/u_add_PartRem_2_39/n2 ), 
        .Y(\u_div/CryTmp[39][6] ) );
  XNOR2X1 U288 ( .A(\u_div/PartRem[40][3] ), .B(\u_div/PartRem[40][2] ), .Y(
        \u_div/SumTmp[39][3] ) );
  OR2X1 U289 ( .A(\u_div/PartRem[39][5] ), .B(\u_div/u_add_PartRem_2_38/n2 ), 
        .Y(\u_div/CryTmp[38][6] ) );
  XNOR2X1 U290 ( .A(\u_div/PartRem[39][3] ), .B(\u_div/PartRem[39][2] ), .Y(
        \u_div/SumTmp[38][3] ) );
  OR2X1 U291 ( .A(\u_div/PartRem[38][5] ), .B(\u_div/u_add_PartRem_2_37/n2 ), 
        .Y(\u_div/CryTmp[37][6] ) );
  XNOR2X1 U292 ( .A(\u_div/PartRem[38][3] ), .B(\u_div/PartRem[38][2] ), .Y(
        \u_div/SumTmp[37][3] ) );
  OR2X1 U293 ( .A(\u_div/PartRem[37][5] ), .B(\u_div/u_add_PartRem_2_36/n2 ), 
        .Y(\u_div/CryTmp[36][6] ) );
  XNOR2X1 U294 ( .A(\u_div/PartRem[37][3] ), .B(\u_div/PartRem[37][2] ), .Y(
        \u_div/SumTmp[36][3] ) );
  OR2X1 U295 ( .A(\u_div/PartRem[36][5] ), .B(\u_div/u_add_PartRem_2_35/n2 ), 
        .Y(\u_div/CryTmp[35][6] ) );
  XNOR2X1 U296 ( .A(\u_div/PartRem[36][3] ), .B(\u_div/PartRem[36][2] ), .Y(
        \u_div/SumTmp[35][3] ) );
  OR2X1 U297 ( .A(\u_div/PartRem[35][5] ), .B(\u_div/u_add_PartRem_2_34/n2 ), 
        .Y(\u_div/CryTmp[34][6] ) );
  XNOR2X1 U298 ( .A(\u_div/PartRem[35][3] ), .B(\u_div/PartRem[35][2] ), .Y(
        \u_div/SumTmp[34][3] ) );
  OR2X1 U299 ( .A(\u_div/PartRem[34][5] ), .B(\u_div/u_add_PartRem_2_33/n2 ), 
        .Y(\u_div/CryTmp[33][6] ) );
  XNOR2X1 U300 ( .A(\u_div/PartRem[34][3] ), .B(\u_div/PartRem[34][2] ), .Y(
        \u_div/SumTmp[33][3] ) );
  OR2X1 U301 ( .A(\u_div/PartRem[33][5] ), .B(\u_div/u_add_PartRem_2_32/n2 ), 
        .Y(\u_div/CryTmp[32][6] ) );
  XNOR2X1 U302 ( .A(\u_div/PartRem[33][3] ), .B(\u_div/PartRem[33][2] ), .Y(
        \u_div/SumTmp[32][3] ) );
  OR2X1 U303 ( .A(\u_div/PartRem[32][5] ), .B(\u_div/u_add_PartRem_2_31/n2 ), 
        .Y(\u_div/CryTmp[31][6] ) );
  XNOR2X1 U304 ( .A(\u_div/PartRem[32][3] ), .B(\u_div/PartRem[32][2] ), .Y(
        \u_div/SumTmp[31][3] ) );
  OR2X1 U305 ( .A(\u_div/PartRem[31][5] ), .B(\u_div/u_add_PartRem_2_30/n2 ), 
        .Y(\u_div/CryTmp[30][6] ) );
  XNOR2X1 U306 ( .A(\u_div/PartRem[31][3] ), .B(\u_div/PartRem[31][2] ), .Y(
        \u_div/SumTmp[30][3] ) );
  OR2X1 U307 ( .A(\u_div/PartRem[30][5] ), .B(\u_div/u_add_PartRem_2_29/n2 ), 
        .Y(\u_div/CryTmp[29][6] ) );
  XNOR2X1 U308 ( .A(\u_div/PartRem[30][3] ), .B(\u_div/PartRem[30][2] ), .Y(
        \u_div/SumTmp[29][3] ) );
  OR2X1 U309 ( .A(\u_div/PartRem[29][5] ), .B(\u_div/u_add_PartRem_2_28/n2 ), 
        .Y(\u_div/CryTmp[28][6] ) );
  XNOR2X1 U310 ( .A(\u_div/PartRem[29][3] ), .B(\u_div/PartRem[29][2] ), .Y(
        \u_div/SumTmp[28][3] ) );
  OR2X1 U311 ( .A(\u_div/PartRem[28][5] ), .B(\u_div/u_add_PartRem_2_27/n2 ), 
        .Y(\u_div/CryTmp[27][6] ) );
  XNOR2X1 U312 ( .A(\u_div/PartRem[28][3] ), .B(\u_div/PartRem[28][2] ), .Y(
        \u_div/SumTmp[27][3] ) );
  OR2X1 U313 ( .A(\u_div/PartRem[27][5] ), .B(\u_div/u_add_PartRem_2_26/n2 ), 
        .Y(\u_div/CryTmp[26][6] ) );
  XNOR2X1 U314 ( .A(\u_div/PartRem[27][3] ), .B(\u_div/PartRem[27][2] ), .Y(
        \u_div/SumTmp[26][3] ) );
  OR2X1 U315 ( .A(\u_div/PartRem[26][5] ), .B(\u_div/u_add_PartRem_2_25/n2 ), 
        .Y(\u_div/CryTmp[25][6] ) );
  XNOR2X1 U316 ( .A(\u_div/PartRem[26][3] ), .B(\u_div/PartRem[26][2] ), .Y(
        \u_div/SumTmp[25][3] ) );
  OR2X1 U317 ( .A(\u_div/PartRem[25][5] ), .B(\u_div/u_add_PartRem_2_24/n2 ), 
        .Y(\u_div/CryTmp[24][6] ) );
  XNOR2X1 U318 ( .A(\u_div/PartRem[25][3] ), .B(\u_div/PartRem[25][2] ), .Y(
        \u_div/SumTmp[24][3] ) );
  OR2X1 U319 ( .A(\u_div/PartRem[24][5] ), .B(\u_div/u_add_PartRem_2_23/n2 ), 
        .Y(\u_div/CryTmp[23][6] ) );
  XNOR2X1 U320 ( .A(\u_div/PartRem[24][3] ), .B(\u_div/PartRem[24][2] ), .Y(
        \u_div/SumTmp[23][3] ) );
  OR2X1 U321 ( .A(\u_div/PartRem[23][5] ), .B(\u_div/u_add_PartRem_2_22/n2 ), 
        .Y(\u_div/CryTmp[22][6] ) );
  XNOR2X1 U322 ( .A(\u_div/PartRem[23][3] ), .B(\u_div/PartRem[23][2] ), .Y(
        \u_div/SumTmp[22][3] ) );
  OR2X1 U323 ( .A(\u_div/PartRem[22][5] ), .B(\u_div/u_add_PartRem_2_21/n2 ), 
        .Y(\u_div/CryTmp[21][6] ) );
  XNOR2X1 U324 ( .A(\u_div/PartRem[22][3] ), .B(\u_div/PartRem[22][2] ), .Y(
        \u_div/SumTmp[21][3] ) );
  OR2X1 U325 ( .A(\u_div/PartRem[21][5] ), .B(\u_div/u_add_PartRem_2_20/n2 ), 
        .Y(\u_div/CryTmp[20][6] ) );
  XNOR2X1 U326 ( .A(\u_div/PartRem[21][3] ), .B(\u_div/PartRem[21][2] ), .Y(
        \u_div/SumTmp[20][3] ) );
  OR2X1 U327 ( .A(\u_div/PartRem[20][5] ), .B(\u_div/u_add_PartRem_2_19/n2 ), 
        .Y(\u_div/CryTmp[19][6] ) );
  XNOR2X1 U328 ( .A(\u_div/PartRem[20][3] ), .B(\u_div/PartRem[20][2] ), .Y(
        \u_div/SumTmp[19][3] ) );
  OR2X1 U329 ( .A(\u_div/PartRem[19][5] ), .B(\u_div/u_add_PartRem_2_18/n2 ), 
        .Y(\u_div/CryTmp[18][6] ) );
  XNOR2X1 U330 ( .A(\u_div/PartRem[19][3] ), .B(\u_div/PartRem[19][2] ), .Y(
        \u_div/SumTmp[18][3] ) );
  OR2X1 U331 ( .A(\u_div/PartRem[18][5] ), .B(\u_div/u_add_PartRem_2_17/n2 ), 
        .Y(\u_div/CryTmp[17][6] ) );
  XNOR2X1 U332 ( .A(\u_div/PartRem[18][3] ), .B(\u_div/PartRem[18][2] ), .Y(
        \u_div/SumTmp[17][3] ) );
  XNOR2X1 U333 ( .A(\u_div/PartRem[17][3] ), .B(\u_div/PartRem[17][2] ), .Y(
        \u_div/SumTmp[16][3] ) );
  OR2X1 U334 ( .A(\u_div/PartRem[16][5] ), .B(\u_div/u_add_PartRem_2_15/n2 ), 
        .Y(\u_div/CryTmp[15][6] ) );
  XNOR2X1 U335 ( .A(\u_div/PartRem[16][3] ), .B(\u_div/PartRem[16][2] ), .Y(
        \u_div/SumTmp[15][3] ) );
  OR2X1 U336 ( .A(\u_div/PartRem[15][5] ), .B(\u_div/u_add_PartRem_2_14/n2 ), 
        .Y(\u_div/CryTmp[14][6] ) );
  XNOR2X1 U337 ( .A(\u_div/PartRem[15][3] ), .B(\u_div/PartRem[15][2] ), .Y(
        \u_div/SumTmp[14][3] ) );
  OR2X1 U338 ( .A(\u_div/PartRem[14][5] ), .B(\u_div/u_add_PartRem_2_13/n2 ), 
        .Y(\u_div/CryTmp[13][6] ) );
  XNOR2X1 U339 ( .A(\u_div/PartRem[14][3] ), .B(\u_div/PartRem[14][2] ), .Y(
        \u_div/SumTmp[13][3] ) );
  OR2X1 U340 ( .A(\u_div/PartRem[13][5] ), .B(\u_div/u_add_PartRem_2_12/n2 ), 
        .Y(\u_div/CryTmp[12][6] ) );
  XNOR2X1 U341 ( .A(\u_div/PartRem[13][3] ), .B(\u_div/PartRem[13][2] ), .Y(
        \u_div/SumTmp[12][3] ) );
  XNOR2X1 U342 ( .A(\u_div/PartRem[12][3] ), .B(\u_div/PartRem[12][2] ), .Y(
        \u_div/SumTmp[11][3] ) );
  OR2X1 U343 ( .A(\u_div/PartRem[11][5] ), .B(\u_div/u_add_PartRem_2_10/n2 ), 
        .Y(\u_div/CryTmp[10][6] ) );
  XNOR2X1 U344 ( .A(\u_div/PartRem[11][3] ), .B(\u_div/PartRem[11][2] ), .Y(
        \u_div/SumTmp[10][3] ) );
  OR2X1 U345 ( .A(\u_div/PartRem[10][5] ), .B(\u_div/u_add_PartRem_2_9/n2 ), 
        .Y(\u_div/CryTmp[9][6] ) );
  XNOR2X1 U346 ( .A(\u_div/PartRem[10][3] ), .B(\u_div/PartRem[10][2] ), .Y(
        \u_div/SumTmp[9][3] ) );
  OR2X1 U347 ( .A(\u_div/PartRem[9][5] ), .B(\u_div/u_add_PartRem_2_8/n2 ), 
        .Y(\u_div/CryTmp[8][6] ) );
  XNOR2X1 U348 ( .A(\u_div/PartRem[9][3] ), .B(\u_div/PartRem[9][2] ), .Y(
        \u_div/SumTmp[8][3] ) );
  OR2X1 U349 ( .A(\u_div/PartRem[8][5] ), .B(\u_div/u_add_PartRem_2_7/n2 ), 
        .Y(\u_div/CryTmp[7][6] ) );
  XNOR2X1 U350 ( .A(\u_div/PartRem[8][3] ), .B(\u_div/PartRem[8][2] ), .Y(
        \u_div/SumTmp[7][3] ) );
  OR2X1 U351 ( .A(\u_div/PartRem[7][5] ), .B(\u_div/u_add_PartRem_2_6/n2 ), 
        .Y(\u_div/CryTmp[6][6] ) );
  XNOR2X1 U352 ( .A(\u_div/PartRem[7][3] ), .B(\u_div/PartRem[7][2] ), .Y(
        \u_div/SumTmp[6][3] ) );
  OR2X1 U353 ( .A(\u_div/PartRem[6][5] ), .B(\u_div/u_add_PartRem_2_5/n2 ), 
        .Y(\u_div/CryTmp[5][6] ) );
  XNOR2X1 U354 ( .A(\u_div/PartRem[6][3] ), .B(\u_div/PartRem[6][2] ), .Y(
        \u_div/SumTmp[5][3] ) );
  OR2X1 U355 ( .A(\u_div/PartRem[5][5] ), .B(\u_div/u_add_PartRem_2_4/n2 ), 
        .Y(\u_div/CryTmp[4][6] ) );
  XNOR2X1 U356 ( .A(\u_div/PartRem[5][3] ), .B(\u_div/PartRem[5][2] ), .Y(
        \u_div/SumTmp[4][3] ) );
  XNOR2X1 U357 ( .A(\u_div/PartRem[4][3] ), .B(\u_div/PartRem[4][2] ), .Y(
        \u_div/SumTmp[3][3] ) );
  XNOR2X1 U358 ( .A(\u_div/PartRem[3][3] ), .B(\u_div/PartRem[3][2] ), .Y(
        \u_div/SumTmp[2][3] ) );
  OR2X1 U359 ( .A(\u_div/PartRem[3][2] ), .B(\u_div/PartRem[3][3] ), .Y(
        \u_div/u_add_PartRem_2_2/n3 ) );
  XNOR2X1 U360 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/PartRem[2][2] ), .Y(
        \u_div/SumTmp[1][3] ) );
  XNOR2X1 U361 ( .A(\u_div/PartRem[63][0] ), .B(\u_div/PartRem[62][0] ), .Y(
        \u_div/SumTmp[59][3] ) );
  XOR2X1 U362 ( .A(\u_div/CryTmp[9][6] ), .B(n2), .Y(\u_div/QInv[9] ) );
  XOR2X1 U363 ( .A(\u_div/CryTmp[8][6] ), .B(n2), .Y(\u_div/QInv[8] ) );
  XOR2X1 U364 ( .A(\u_div/CryTmp[5][6] ), .B(n3), .Y(\u_div/QInv[5] ) );
  XOR2X1 U365 ( .A(\u_div/CryTmp[59][6] ), .B(n2), .Y(\u_div/QInv[59] ) );
  XOR2X1 U366 ( .A(\u_div/CryTmp[58][6] ), .B(n4), .Y(\u_div/QInv[58] ) );
  XOR2X1 U367 ( .A(\u_div/CryTmp[57][6] ), .B(n3), .Y(\u_div/QInv[57] ) );
  XOR2X1 U368 ( .A(\u_div/CryTmp[56][6] ), .B(n2), .Y(\u_div/QInv[56] ) );
  XOR2X1 U369 ( .A(\u_div/CryTmp[55][6] ), .B(n4), .Y(\u_div/QInv[55] ) );
  XOR2X1 U370 ( .A(\u_div/CryTmp[54][6] ), .B(n3), .Y(\u_div/QInv[54] ) );
  XOR2X1 U371 ( .A(\u_div/CryTmp[52][6] ), .B(n4), .Y(\u_div/QInv[52] ) );
  XOR2X1 U372 ( .A(\u_div/CryTmp[51][6] ), .B(n3), .Y(\u_div/QInv[51] ) );
  XOR2X1 U373 ( .A(\u_div/CryTmp[50][6] ), .B(n2), .Y(\u_div/QInv[50] ) );
  XOR2X1 U374 ( .A(\u_div/CryTmp[4][6] ), .B(n4), .Y(\u_div/QInv[4] ) );
  XOR2X1 U375 ( .A(\u_div/CryTmp[49][6] ), .B(n3), .Y(\u_div/QInv[49] ) );
  XOR2X1 U376 ( .A(\u_div/CryTmp[44][6] ), .B(n4), .Y(\u_div/QInv[44] ) );
  XOR2X1 U377 ( .A(\u_div/CryTmp[43][6] ), .B(n3), .Y(\u_div/QInv[43] ) );
  XOR2X1 U378 ( .A(\u_div/CryTmp[42][6] ), .B(n2), .Y(\u_div/QInv[42] ) );
  XOR2X1 U379 ( .A(\u_div/CryTmp[41][6] ), .B(n4), .Y(\u_div/QInv[41] ) );
  XOR2X1 U380 ( .A(\u_div/CryTmp[40][6] ), .B(n3), .Y(\u_div/QInv[40] ) );
  XOR2X1 U381 ( .A(\u_div/CryTmp[3][6] ), .B(n2), .Y(\u_div/QInv[3] ) );
  XOR2X1 U382 ( .A(\u_div/CryTmp[39][6] ), .B(n4), .Y(\u_div/QInv[39] ) );
  XOR2X1 U383 ( .A(\u_div/CryTmp[38][6] ), .B(n3), .Y(\u_div/QInv[38] ) );
  XOR2X1 U384 ( .A(\u_div/CryTmp[37][6] ), .B(n2), .Y(\u_div/QInv[37] ) );
  XOR2X1 U385 ( .A(\u_div/CryTmp[34][6] ), .B(n4), .Y(\u_div/QInv[34] ) );
  XOR2X1 U386 ( .A(\u_div/CryTmp[33][6] ), .B(n3), .Y(\u_div/QInv[33] ) );
  XOR2X1 U387 ( .A(\u_div/CryTmp[32][6] ), .B(n2), .Y(\u_div/QInv[32] ) );
  XOR2X1 U388 ( .A(\u_div/CryTmp[31][6] ), .B(n4), .Y(\u_div/QInv[31] ) );
  XOR2X1 U389 ( .A(\u_div/CryTmp[30][6] ), .B(n3), .Y(\u_div/QInv[30] ) );
  XOR2X1 U390 ( .A(\u_div/CryTmp[2][6] ), .B(n2), .Y(\u_div/QInv[2] ) );
  XOR2X1 U391 ( .A(\u_div/CryTmp[29][6] ), .B(n4), .Y(\u_div/QInv[29] ) );
  XOR2X1 U392 ( .A(\u_div/CryTmp[27][6] ), .B(n2), .Y(\u_div/QInv[27] ) );
  XOR2X1 U393 ( .A(\u_div/CryTmp[26][6] ), .B(n4), .Y(\u_div/QInv[26] ) );
  XOR2X1 U394 ( .A(\u_div/CryTmp[24][6] ), .B(n2), .Y(\u_div/QInv[24] ) );
  XOR2X1 U395 ( .A(\u_div/CryTmp[23][6] ), .B(n4), .Y(\u_div/QInv[23] ) );
  XOR2X1 U396 ( .A(\u_div/CryTmp[22][6] ), .B(n3), .Y(\u_div/QInv[22] ) );
  XOR2X1 U397 ( .A(\u_div/CryTmp[21][6] ), .B(n2), .Y(\u_div/QInv[21] ) );
  XOR2X1 U398 ( .A(\u_div/CryTmp[20][6] ), .B(n4), .Y(\u_div/QInv[20] ) );
  XOR2X1 U399 ( .A(\u_div/CryTmp[1][6] ), .B(n3), .Y(\u_div/QInv[1] ) );
  XOR2X1 U400 ( .A(\u_div/CryTmp[19][6] ), .B(n2), .Y(\u_div/QInv[19] ) );
  XOR2X1 U401 ( .A(\u_div/CryTmp[18][6] ), .B(n4), .Y(\u_div/QInv[18] ) );
  XOR2X1 U402 ( .A(\u_div/CryTmp[16][6] ), .B(n4), .Y(\u_div/QInv[16] ) );
  XOR2X1 U403 ( .A(\u_div/CryTmp[15][6] ), .B(n3), .Y(\u_div/QInv[15] ) );
  XOR2X1 U404 ( .A(\u_div/CryTmp[14][6] ), .B(n4), .Y(\u_div/QInv[14] ) );
  XOR2X1 U405 ( .A(\u_div/CryTmp[13][6] ), .B(n3), .Y(\u_div/QInv[13] ) );
  XOR2X1 U406 ( .A(\u_div/CryTmp[12][6] ), .B(n4), .Y(\u_div/QInv[12] ) );
  XOR2X1 U407 ( .A(\u_div/CryTmp[11][6] ), .B(n3), .Y(\u_div/QInv[11] ) );
  XOR2X1 U408 ( .A(\u_div/CryTmp[10][6] ), .B(n4), .Y(\u_div/QInv[10] ) );
endmodule


module GSIM_DW01_inc_8 ( A, SUM );
  input [63:0] A;
  output [63:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;

  NOR2BX1 U2 ( .AN(A[62]), .B(n21), .Y(n20) );
  NAND2XL U3 ( .A(A[60]), .B(n22), .Y(n23) );
  XOR2X4 U4 ( .A(A[63]), .B(n20), .Y(SUM[63]) );
  NAND3X1 U5 ( .A(A[60]), .B(n22), .C(A[61]), .Y(n21) );
  NOR3BX1 U6 ( .AN(A[55]), .B(n2), .C(n30), .Y(n28) );
  NOR3BX1 U7 ( .AN(A[51]), .B(n3), .C(n34), .Y(n32) );
  NOR3BX1 U8 ( .AN(A[47]), .B(n4), .C(n38), .Y(n36) );
  NOR3BX1 U9 ( .AN(A[43]), .B(n5), .C(n42), .Y(n40) );
  NOR3BX1 U10 ( .AN(A[39]), .B(n6), .C(n46), .Y(n44) );
  NOR3BX1 U11 ( .AN(A[35]), .B(n7), .C(n52), .Y(n50) );
  NOR3BX1 U12 ( .AN(A[31]), .B(n8), .C(n56), .Y(n54) );
  NOR3BX1 U13 ( .AN(A[27]), .B(n9), .C(n60), .Y(n58) );
  NOR3BX1 U14 ( .AN(A[23]), .B(n10), .C(n64), .Y(n62) );
  NOR3BX1 U15 ( .AN(A[19]), .B(n11), .C(n68), .Y(n66) );
  NOR3BX1 U16 ( .AN(A[15]), .B(n12), .C(n72), .Y(n70) );
  NOR3BX1 U17 ( .AN(A[11]), .B(n13), .C(n76), .Y(n74) );
  NOR3BX1 U18 ( .AN(A[7]), .B(n14), .C(n19), .Y(n17) );
  CLKINVX1 U19 ( .A(A[58]), .Y(n1) );
  CLKINVX1 U20 ( .A(A[54]), .Y(n2) );
  CLKINVX1 U21 ( .A(A[50]), .Y(n3) );
  CLKINVX1 U22 ( .A(A[46]), .Y(n4) );
  CLKINVX1 U23 ( .A(A[42]), .Y(n5) );
  CLKINVX1 U24 ( .A(A[38]), .Y(n6) );
  CLKINVX1 U25 ( .A(A[34]), .Y(n7) );
  CLKINVX1 U26 ( .A(A[30]), .Y(n8) );
  CLKINVX1 U27 ( .A(A[26]), .Y(n9) );
  CLKINVX1 U28 ( .A(A[22]), .Y(n10) );
  CLKINVX1 U29 ( .A(A[18]), .Y(n11) );
  CLKINVX1 U30 ( .A(A[14]), .Y(n12) );
  CLKINVX1 U31 ( .A(A[10]), .Y(n13) );
  NAND3X1 U32 ( .A(A[4]), .B(n26), .C(A[5]), .Y(n19) );
  CLKINVX1 U33 ( .A(A[6]), .Y(n14) );
  NOR3BX1 U34 ( .AN(A[3]), .B(n15), .C(n48), .Y(n26) );
  NOR2XL U35 ( .A(n24), .B(n1), .Y(n27) );
  NAND2XL U36 ( .A(A[56]), .B(n28), .Y(n29) );
  NOR2XL U37 ( .A(n30), .B(n2), .Y(n31) );
  NAND2XL U38 ( .A(A[52]), .B(n32), .Y(n33) );
  NOR2XL U39 ( .A(n34), .B(n3), .Y(n35) );
  NAND2XL U40 ( .A(A[48]), .B(n36), .Y(n37) );
  NOR2XL U41 ( .A(n38), .B(n4), .Y(n39) );
  NAND2XL U42 ( .A(A[44]), .B(n40), .Y(n41) );
  NOR2XL U43 ( .A(n42), .B(n5), .Y(n43) );
  NAND2XL U44 ( .A(A[40]), .B(n44), .Y(n45) );
  NOR2XL U45 ( .A(n46), .B(n6), .Y(n49) );
  NAND2XL U46 ( .A(A[36]), .B(n50), .Y(n51) );
  NOR2XL U47 ( .A(n52), .B(n7), .Y(n53) );
  NAND2XL U48 ( .A(A[32]), .B(n54), .Y(n55) );
  NOR2XL U49 ( .A(n56), .B(n8), .Y(n57) );
  NAND2XL U50 ( .A(A[28]), .B(n58), .Y(n59) );
  NOR2XL U51 ( .A(n60), .B(n9), .Y(n61) );
  NAND2XL U52 ( .A(A[24]), .B(n62), .Y(n63) );
  NOR2XL U53 ( .A(n64), .B(n10), .Y(n65) );
  NAND2XL U54 ( .A(A[20]), .B(n66), .Y(n67) );
  NOR2XL U55 ( .A(n68), .B(n11), .Y(n69) );
  NAND2XL U56 ( .A(A[16]), .B(n70), .Y(n71) );
  NOR2XL U57 ( .A(n72), .B(n12), .Y(n73) );
  NAND2XL U58 ( .A(A[12]), .B(n74), .Y(n75) );
  NOR2XL U59 ( .A(n76), .B(n13), .Y(n77) );
  NAND2XL U60 ( .A(A[8]), .B(n17), .Y(n16) );
  NOR2XL U61 ( .A(n19), .B(n14), .Y(n18) );
  NAND2XL U62 ( .A(A[4]), .B(n26), .Y(n25) );
  XOR2XL U63 ( .A(A[60]), .B(n22), .Y(SUM[60]) );
  NOR2XL U64 ( .A(n48), .B(n15), .Y(n47) );
  NOR3BX1 U65 ( .AN(A[59]), .B(n1), .C(n24), .Y(n22) );
  CLKINVX1 U66 ( .A(A[2]), .Y(n15) );
  XNOR2X1 U67 ( .A(A[9]), .B(n16), .Y(SUM[9]) );
  XOR2X1 U68 ( .A(A[8]), .B(n17), .Y(SUM[8]) );
  XOR2X1 U69 ( .A(A[7]), .B(n18), .Y(SUM[7]) );
  XOR2X1 U70 ( .A(n14), .B(n19), .Y(SUM[6]) );
  XNOR2X1 U71 ( .A(A[62]), .B(n21), .Y(SUM[62]) );
  XNOR2X1 U72 ( .A(A[61]), .B(n23), .Y(SUM[61]) );
  XNOR2X1 U73 ( .A(A[5]), .B(n25), .Y(SUM[5]) );
  XOR2X1 U74 ( .A(A[59]), .B(n27), .Y(SUM[59]) );
  XOR2X1 U75 ( .A(n1), .B(n24), .Y(SUM[58]) );
  NAND3X1 U76 ( .A(A[56]), .B(n28), .C(A[57]), .Y(n24) );
  XNOR2X1 U77 ( .A(A[57]), .B(n29), .Y(SUM[57]) );
  XOR2X1 U78 ( .A(A[56]), .B(n28), .Y(SUM[56]) );
  XOR2X1 U79 ( .A(A[55]), .B(n31), .Y(SUM[55]) );
  XOR2X1 U80 ( .A(n2), .B(n30), .Y(SUM[54]) );
  NAND3X1 U81 ( .A(A[52]), .B(n32), .C(A[53]), .Y(n30) );
  XNOR2X1 U82 ( .A(A[53]), .B(n33), .Y(SUM[53]) );
  XOR2X1 U83 ( .A(A[52]), .B(n32), .Y(SUM[52]) );
  XOR2X1 U84 ( .A(A[51]), .B(n35), .Y(SUM[51]) );
  XOR2X1 U85 ( .A(n3), .B(n34), .Y(SUM[50]) );
  NAND3X1 U86 ( .A(A[48]), .B(n36), .C(A[49]), .Y(n34) );
  XOR2X1 U87 ( .A(A[4]), .B(n26), .Y(SUM[4]) );
  XNOR2X1 U88 ( .A(A[49]), .B(n37), .Y(SUM[49]) );
  XOR2X1 U89 ( .A(A[48]), .B(n36), .Y(SUM[48]) );
  XOR2X1 U90 ( .A(A[47]), .B(n39), .Y(SUM[47]) );
  XOR2X1 U91 ( .A(n4), .B(n38), .Y(SUM[46]) );
  NAND3X1 U92 ( .A(A[44]), .B(n40), .C(A[45]), .Y(n38) );
  XNOR2X1 U93 ( .A(A[45]), .B(n41), .Y(SUM[45]) );
  XOR2X1 U94 ( .A(A[44]), .B(n40), .Y(SUM[44]) );
  XOR2X1 U95 ( .A(A[43]), .B(n43), .Y(SUM[43]) );
  XOR2X1 U96 ( .A(n5), .B(n42), .Y(SUM[42]) );
  NAND3X1 U97 ( .A(A[40]), .B(n44), .C(A[41]), .Y(n42) );
  XNOR2X1 U98 ( .A(A[41]), .B(n45), .Y(SUM[41]) );
  XOR2X1 U99 ( .A(A[40]), .B(n44), .Y(SUM[40]) );
  XOR2X1 U100 ( .A(A[3]), .B(n47), .Y(SUM[3]) );
  XOR2X1 U101 ( .A(A[39]), .B(n49), .Y(SUM[39]) );
  XOR2X1 U102 ( .A(n6), .B(n46), .Y(SUM[38]) );
  NAND3X1 U103 ( .A(A[36]), .B(n50), .C(A[37]), .Y(n46) );
  XNOR2X1 U104 ( .A(A[37]), .B(n51), .Y(SUM[37]) );
  XOR2X1 U105 ( .A(A[36]), .B(n50), .Y(SUM[36]) );
  XOR2X1 U106 ( .A(A[35]), .B(n53), .Y(SUM[35]) );
  XOR2X1 U107 ( .A(n7), .B(n52), .Y(SUM[34]) );
  NAND3X1 U108 ( .A(A[32]), .B(n54), .C(A[33]), .Y(n52) );
  XNOR2X1 U109 ( .A(A[33]), .B(n55), .Y(SUM[33]) );
  XOR2X1 U110 ( .A(A[32]), .B(n54), .Y(SUM[32]) );
  XOR2X1 U111 ( .A(A[31]), .B(n57), .Y(SUM[31]) );
  XOR2X1 U112 ( .A(n8), .B(n56), .Y(SUM[30]) );
  NAND3X1 U113 ( .A(A[28]), .B(n58), .C(A[29]), .Y(n56) );
  XOR2X1 U114 ( .A(n15), .B(n48), .Y(SUM[2]) );
  XNOR2X1 U115 ( .A(A[29]), .B(n59), .Y(SUM[29]) );
  XOR2X1 U116 ( .A(A[28]), .B(n58), .Y(SUM[28]) );
  XOR2X1 U117 ( .A(A[27]), .B(n61), .Y(SUM[27]) );
  XOR2X1 U118 ( .A(n9), .B(n60), .Y(SUM[26]) );
  NAND3X1 U119 ( .A(A[24]), .B(n62), .C(A[25]), .Y(n60) );
  XNOR2X1 U120 ( .A(A[25]), .B(n63), .Y(SUM[25]) );
  XOR2X1 U121 ( .A(A[24]), .B(n62), .Y(SUM[24]) );
  XOR2X1 U122 ( .A(A[23]), .B(n65), .Y(SUM[23]) );
  XOR2X1 U123 ( .A(n10), .B(n64), .Y(SUM[22]) );
  NAND3X1 U124 ( .A(A[20]), .B(n66), .C(A[21]), .Y(n64) );
  XNOR2X1 U125 ( .A(A[21]), .B(n67), .Y(SUM[21]) );
  XOR2X1 U126 ( .A(A[20]), .B(n66), .Y(SUM[20]) );
  XOR2X1 U127 ( .A(A[19]), .B(n69), .Y(SUM[19]) );
  XOR2X1 U128 ( .A(n11), .B(n68), .Y(SUM[18]) );
  NAND3X1 U129 ( .A(A[16]), .B(n70), .C(A[17]), .Y(n68) );
  XNOR2X1 U130 ( .A(A[17]), .B(n71), .Y(SUM[17]) );
  XOR2X1 U131 ( .A(A[16]), .B(n70), .Y(SUM[16]) );
  XOR2X1 U132 ( .A(A[15]), .B(n73), .Y(SUM[15]) );
  XOR2X1 U133 ( .A(n12), .B(n72), .Y(SUM[14]) );
  NAND3X1 U134 ( .A(A[12]), .B(n74), .C(A[13]), .Y(n72) );
  XNOR2X1 U135 ( .A(A[13]), .B(n75), .Y(SUM[13]) );
  XOR2X1 U136 ( .A(A[12]), .B(n74), .Y(SUM[12]) );
  XOR2X1 U137 ( .A(A[11]), .B(n77), .Y(SUM[11]) );
  XOR2X1 U138 ( .A(n13), .B(n76), .Y(SUM[10]) );
  NAND3X1 U139 ( .A(A[8]), .B(n17), .C(A[9]), .Y(n76) );
  NAND2X1 U140 ( .A(A[1]), .B(A[0]), .Y(n48) );
endmodule


module GSIM_DW01_absval_6 ( A, ABSVAL );
  input [63:0] A;
  output [63:0] ABSVAL;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69;
  wire   [63:0] AMUX1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  GSIM_DW01_inc_8 NEG ( .A({n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
        n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
        n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
        n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, 
        n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69}), .SUM({
        AMUX1[63:2], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1}) );
  CLKMX2X2 U1 ( .A(A[61]), .B(AMUX1[61]), .S0(n4), .Y(ABSVAL[61]) );
  CLKINVX1 U2 ( .A(A[60]), .Y(n9) );
  CLKINVX1 U3 ( .A(A[58]), .Y(n11) );
  CLKINVX1 U4 ( .A(A[56]), .Y(n13) );
  CLKINVX1 U5 ( .A(A[52]), .Y(n17) );
  CLKINVX1 U6 ( .A(A[54]), .Y(n15) );
  CLKINVX1 U7 ( .A(A[50]), .Y(n19) );
  CLKINVX1 U8 ( .A(A[48]), .Y(n21) );
  CLKINVX1 U9 ( .A(A[46]), .Y(n23) );
  CLKINVX1 U10 ( .A(A[44]), .Y(n25) );
  CLKINVX1 U11 ( .A(A[40]), .Y(n29) );
  CLKINVX1 U12 ( .A(A[42]), .Y(n27) );
  CLKINVX1 U13 ( .A(A[38]), .Y(n31) );
  CLKINVX1 U14 ( .A(A[36]), .Y(n33) );
  CLKINVX1 U15 ( .A(A[34]), .Y(n35) );
  CLKINVX1 U16 ( .A(A[32]), .Y(n37) );
  CLKINVX1 U17 ( .A(A[28]), .Y(n41) );
  CLKINVX1 U18 ( .A(A[30]), .Y(n39) );
  CLKINVX1 U19 ( .A(A[26]), .Y(n43) );
  CLKINVX1 U20 ( .A(A[24]), .Y(n45) );
  CLKINVX1 U21 ( .A(A[22]), .Y(n47) );
  CLKINVX1 U22 ( .A(A[20]), .Y(n49) );
  CLKINVX1 U23 ( .A(A[16]), .Y(n53) );
  CLKINVX1 U24 ( .A(A[18]), .Y(n51) );
  CLKINVX1 U25 ( .A(A[14]), .Y(n55) );
  CLKINVX1 U26 ( .A(A[12]), .Y(n57) );
  CLKINVX1 U27 ( .A(A[6]), .Y(n63) );
  CLKINVX1 U28 ( .A(A[8]), .Y(n61) );
  CLKINVX1 U29 ( .A(A[10]), .Y(n59) );
  CLKBUFX2 U30 ( .A(n6), .Y(n5) );
  INVX3 U31 ( .A(n6), .Y(n4) );
  INVX3 U32 ( .A(n5), .Y(n3) );
  INVX3 U33 ( .A(n5), .Y(n2) );
  INVX3 U34 ( .A(n5), .Y(n1) );
  CLKINVX1 U35 ( .A(A[63]), .Y(n6) );
  CLKINVX1 U36 ( .A(A[3]), .Y(n66) );
  CLKINVX1 U37 ( .A(A[2]), .Y(n67) );
  CLKINVX1 U38 ( .A(A[5]), .Y(n64) );
  CLKINVX1 U39 ( .A(A[62]), .Y(n7) );
  CLKINVX1 U40 ( .A(A[15]), .Y(n54) );
  CLKINVX1 U41 ( .A(A[11]), .Y(n58) );
  CLKINVX1 U42 ( .A(A[7]), .Y(n62) );
  CLKINVX1 U43 ( .A(A[4]), .Y(n65) );
  CLKINVX1 U44 ( .A(A[59]), .Y(n10) );
  CLKINVX1 U45 ( .A(A[45]), .Y(n24) );
  CLKINVX1 U46 ( .A(A[33]), .Y(n36) );
  CLKINVX1 U47 ( .A(A[29]), .Y(n40) );
  CLKINVX1 U48 ( .A(A[25]), .Y(n44) );
  CLKINVX1 U49 ( .A(A[21]), .Y(n48) );
  CLKINVX1 U50 ( .A(A[17]), .Y(n52) );
  CLKINVX1 U51 ( .A(A[13]), .Y(n56) );
  CLKINVX1 U52 ( .A(A[9]), .Y(n60) );
  CLKINVX1 U53 ( .A(A[55]), .Y(n14) );
  CLKINVX1 U54 ( .A(A[51]), .Y(n18) );
  CLKINVX1 U55 ( .A(A[47]), .Y(n22) );
  CLKINVX1 U56 ( .A(A[43]), .Y(n26) );
  CLKINVX1 U57 ( .A(A[39]), .Y(n30) );
  CLKINVX1 U58 ( .A(A[35]), .Y(n34) );
  CLKINVX1 U59 ( .A(A[31]), .Y(n38) );
  CLKINVX1 U60 ( .A(A[27]), .Y(n42) );
  CLKINVX1 U61 ( .A(A[23]), .Y(n46) );
  CLKINVX1 U62 ( .A(A[19]), .Y(n50) );
  CLKINVX1 U63 ( .A(A[57]), .Y(n12) );
  CLKINVX1 U64 ( .A(A[53]), .Y(n16) );
  CLKINVX1 U65 ( .A(A[49]), .Y(n20) );
  CLKINVX1 U66 ( .A(A[41]), .Y(n28) );
  CLKINVX1 U67 ( .A(A[37]), .Y(n32) );
  CLKINVX1 U68 ( .A(A[0]), .Y(n69) );
  CLKINVX1 U69 ( .A(A[1]), .Y(n68) );
  CLKINVX1 U70 ( .A(A[61]), .Y(n8) );
  CLKMX2X2 U71 ( .A(A[9]), .B(AMUX1[9]), .S0(n3), .Y(ABSVAL[9]) );
  CLKMX2X2 U72 ( .A(A[8]), .B(AMUX1[8]), .S0(n4), .Y(ABSVAL[8]) );
  CLKMX2X2 U73 ( .A(A[7]), .B(AMUX1[7]), .S0(n4), .Y(ABSVAL[7]) );
  CLKMX2X2 U74 ( .A(A[6]), .B(AMUX1[6]), .S0(n4), .Y(ABSVAL[6]) );
  AND2X1 U75 ( .A(AMUX1[63]), .B(n4), .Y(ABSVAL[63]) );
  CLKMX2X2 U76 ( .A(A[62]), .B(AMUX1[62]), .S0(n4), .Y(ABSVAL[62]) );
  CLKMX2X2 U77 ( .A(A[60]), .B(AMUX1[60]), .S0(n4), .Y(ABSVAL[60]) );
  CLKMX2X2 U78 ( .A(A[5]), .B(AMUX1[5]), .S0(n4), .Y(ABSVAL[5]) );
  CLKMX2X2 U79 ( .A(A[59]), .B(AMUX1[59]), .S0(n4), .Y(ABSVAL[59]) );
  CLKMX2X2 U80 ( .A(A[58]), .B(AMUX1[58]), .S0(n4), .Y(ABSVAL[58]) );
  CLKMX2X2 U81 ( .A(A[57]), .B(AMUX1[57]), .S0(n4), .Y(ABSVAL[57]) );
  CLKMX2X2 U82 ( .A(A[56]), .B(AMUX1[56]), .S0(n3), .Y(ABSVAL[56]) );
  CLKMX2X2 U83 ( .A(A[55]), .B(AMUX1[55]), .S0(n3), .Y(ABSVAL[55]) );
  CLKMX2X2 U84 ( .A(A[54]), .B(AMUX1[54]), .S0(n3), .Y(ABSVAL[54]) );
  CLKMX2X2 U85 ( .A(A[53]), .B(AMUX1[53]), .S0(n3), .Y(ABSVAL[53]) );
  CLKMX2X2 U86 ( .A(A[52]), .B(AMUX1[52]), .S0(n3), .Y(ABSVAL[52]) );
  CLKMX2X2 U87 ( .A(A[51]), .B(AMUX1[51]), .S0(n3), .Y(ABSVAL[51]) );
  CLKMX2X2 U88 ( .A(A[50]), .B(AMUX1[50]), .S0(n3), .Y(ABSVAL[50]) );
  CLKMX2X2 U89 ( .A(A[4]), .B(AMUX1[4]), .S0(n3), .Y(ABSVAL[4]) );
  CLKMX2X2 U90 ( .A(A[49]), .B(AMUX1[49]), .S0(n3), .Y(ABSVAL[49]) );
  CLKMX2X2 U91 ( .A(A[48]), .B(AMUX1[48]), .S0(n3), .Y(ABSVAL[48]) );
  CLKMX2X2 U92 ( .A(A[47]), .B(AMUX1[47]), .S0(n3), .Y(ABSVAL[47]) );
  CLKMX2X2 U93 ( .A(A[46]), .B(AMUX1[46]), .S0(n3), .Y(ABSVAL[46]) );
  CLKMX2X2 U94 ( .A(A[45]), .B(AMUX1[45]), .S0(n3), .Y(ABSVAL[45]) );
  CLKMX2X2 U95 ( .A(A[44]), .B(AMUX1[44]), .S0(n2), .Y(ABSVAL[44]) );
  CLKMX2X2 U96 ( .A(A[43]), .B(AMUX1[43]), .S0(n2), .Y(ABSVAL[43]) );
  CLKMX2X2 U97 ( .A(A[42]), .B(AMUX1[42]), .S0(n2), .Y(ABSVAL[42]) );
  CLKMX2X2 U98 ( .A(A[41]), .B(AMUX1[41]), .S0(n2), .Y(ABSVAL[41]) );
  CLKMX2X2 U99 ( .A(A[40]), .B(AMUX1[40]), .S0(n2), .Y(ABSVAL[40]) );
  CLKMX2X2 U100 ( .A(A[3]), .B(AMUX1[3]), .S0(n2), .Y(ABSVAL[3]) );
  CLKMX2X2 U101 ( .A(A[39]), .B(AMUX1[39]), .S0(n2), .Y(ABSVAL[39]) );
  CLKMX2X2 U102 ( .A(A[38]), .B(AMUX1[38]), .S0(n2), .Y(ABSVAL[38]) );
  CLKMX2X2 U103 ( .A(A[37]), .B(AMUX1[37]), .S0(n2), .Y(ABSVAL[37]) );
  CLKMX2X2 U104 ( .A(A[36]), .B(AMUX1[36]), .S0(n2), .Y(ABSVAL[36]) );
  CLKMX2X2 U105 ( .A(A[35]), .B(AMUX1[35]), .S0(n2), .Y(ABSVAL[35]) );
  CLKMX2X2 U106 ( .A(A[34]), .B(AMUX1[34]), .S0(n2), .Y(ABSVAL[34]) );
  CLKMX2X2 U107 ( .A(A[33]), .B(AMUX1[33]), .S0(n1), .Y(ABSVAL[33]) );
  CLKMX2X2 U108 ( .A(A[32]), .B(AMUX1[32]), .S0(n1), .Y(ABSVAL[32]) );
  CLKMX2X2 U109 ( .A(A[31]), .B(AMUX1[31]), .S0(n1), .Y(ABSVAL[31]) );
  CLKMX2X2 U110 ( .A(A[30]), .B(AMUX1[30]), .S0(n1), .Y(ABSVAL[30]) );
  CLKMX2X2 U111 ( .A(A[2]), .B(AMUX1[2]), .S0(n1), .Y(ABSVAL[2]) );
  CLKMX2X2 U112 ( .A(A[29]), .B(AMUX1[29]), .S0(n1), .Y(ABSVAL[29]) );
  CLKMX2X2 U113 ( .A(A[28]), .B(AMUX1[28]), .S0(n1), .Y(ABSVAL[28]) );
  CLKMX2X2 U114 ( .A(A[27]), .B(AMUX1[27]), .S0(n1), .Y(ABSVAL[27]) );
  CLKMX2X2 U115 ( .A(A[26]), .B(AMUX1[26]), .S0(n1), .Y(ABSVAL[26]) );
  CLKMX2X2 U116 ( .A(A[25]), .B(AMUX1[25]), .S0(n1), .Y(ABSVAL[25]) );
  CLKMX2X2 U117 ( .A(A[24]), .B(AMUX1[24]), .S0(n1), .Y(ABSVAL[24]) );
  CLKMX2X2 U118 ( .A(A[23]), .B(AMUX1[23]), .S0(n1), .Y(ABSVAL[23]) );
  CLKMX2X2 U119 ( .A(A[22]), .B(AMUX1[22]), .S0(n1), .Y(ABSVAL[22]) );
  CLKMX2X2 U120 ( .A(A[21]), .B(AMUX1[21]), .S0(n1), .Y(ABSVAL[21]) );
  CLKMX2X2 U121 ( .A(A[20]), .B(AMUX1[20]), .S0(n1), .Y(ABSVAL[20]) );
  CLKMX2X2 U122 ( .A(A[19]), .B(AMUX1[19]), .S0(n1), .Y(ABSVAL[19]) );
  CLKMX2X2 U123 ( .A(A[18]), .B(AMUX1[18]), .S0(n1), .Y(ABSVAL[18]) );
  CLKMX2X2 U124 ( .A(A[17]), .B(AMUX1[17]), .S0(n2), .Y(ABSVAL[17]) );
  CLKMX2X2 U125 ( .A(A[16]), .B(AMUX1[16]), .S0(n2), .Y(ABSVAL[16]) );
  CLKMX2X2 U126 ( .A(A[15]), .B(AMUX1[15]), .S0(n2), .Y(ABSVAL[15]) );
  CLKMX2X2 U127 ( .A(A[14]), .B(AMUX1[14]), .S0(n2), .Y(ABSVAL[14]) );
  CLKMX2X2 U128 ( .A(A[13]), .B(AMUX1[13]), .S0(n3), .Y(ABSVAL[13]) );
  CLKMX2X2 U129 ( .A(A[12]), .B(AMUX1[12]), .S0(n3), .Y(ABSVAL[12]) );
  CLKMX2X2 U130 ( .A(A[11]), .B(AMUX1[11]), .S0(n3), .Y(ABSVAL[11]) );
  CLKMX2X2 U131 ( .A(A[10]), .B(AMUX1[10]), .S0(n2), .Y(ABSVAL[10]) );
endmodule


module GSIM_DW_inc_6 ( carry_in, a, carry_out, sum );
  input [63:0] a;
  output [63:0] sum;
  input carry_in;
  output carry_out;
  wire   \sum[63] , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63;
  assign sum[62] = \sum[63] ;
  assign sum[61] = \sum[63] ;
  assign sum[63] = \sum[63] ;

  ADDHXL U12 ( .A(a[54]), .B(n10), .CO(n9), .S(sum[54]) );
  ADDHXL U20 ( .A(a[46]), .B(n18), .CO(n17), .S(sum[46]) );
  ADDHXL U31 ( .A(a[35]), .B(n29), .CO(n28), .S(sum[35]) );
  ADDHXL U41 ( .A(a[25]), .B(n39), .CO(n38), .S(sum[25]) );
  ADDHXL U51 ( .A(a[15]), .B(n49), .CO(n48), .S(sum[15]) );
  ADDHXL U60 ( .A(a[6]), .B(n58), .CO(n57), .S(sum[6]) );
  ADDHXL U70 ( .A(a[53]), .B(n11), .CO(n10), .S(sum[53]) );
  ADDHXL U71 ( .A(a[27]), .B(n37), .CO(n36), .S(sum[27]) );
  ADDHXL U72 ( .A(a[37]), .B(n27), .CO(n26), .S(sum[37]) );
  ADDHXL U73 ( .A(a[26]), .B(n38), .CO(n37), .S(sum[26]) );
  ADDHXL U74 ( .A(a[36]), .B(n28), .CO(n27), .S(sum[36]) );
  ADDHXL U75 ( .A(a[52]), .B(n12), .CO(n11), .S(sum[52]) );
  ADDHX1 U76 ( .A(a[5]), .B(n59), .CO(n58), .S(sum[5]) );
  ADDHX1 U77 ( .A(a[16]), .B(n48), .CO(n47), .S(sum[16]) );
  ADDHX1 U78 ( .A(a[14]), .B(n50), .CO(n49), .S(sum[14]) );
  ADDHX1 U79 ( .A(a[44]), .B(n20), .CO(n19), .S(sum[44]) );
  ADDHX1 U80 ( .A(a[34]), .B(n30), .CO(n29), .S(sum[34]) );
  ADDHX1 U81 ( .A(a[42]), .B(n22), .CO(n21), .S(sum[42]) );
  ADDHX1 U82 ( .A(a[50]), .B(n14), .CO(n13), .S(sum[50]) );
  ADDHX1 U83 ( .A(a[21]), .B(n43), .CO(n42), .S(sum[21]) );
  ADDHX1 U84 ( .A(a[3]), .B(n61), .CO(n60), .S(sum[3]) );
  ADDHX1 U85 ( .A(a[9]), .B(n55), .CO(n54), .S(sum[9]) );
  ADDHX1 U86 ( .A(a[55]), .B(n9), .CO(n8), .S(sum[55]) );
  ADDHX1 U87 ( .A(a[47]), .B(n17), .CO(n16), .S(sum[47]) );
  ADDHX1 U88 ( .A(a[1]), .B(n63), .CO(n62), .S(sum[1]) );
  ADDHX1 U89 ( .A(a[7]), .B(n57), .CO(n56), .S(sum[7]) );
  ADDHX1 U90 ( .A(a[58]), .B(n6), .CO(n5), .S(sum[58]) );
  ADDHX1 U91 ( .A(a[39]), .B(n25), .CO(n24), .S(sum[39]) );
  ADDHX1 U92 ( .A(a[40]), .B(n24), .CO(n23), .S(sum[40]) );
  ADDHX1 U93 ( .A(a[31]), .B(n33), .CO(n32), .S(sum[31]) );
  ADDHX1 U94 ( .A(a[29]), .B(n35), .CO(n34), .S(sum[29]) );
  ADDHX1 U95 ( .A(a[23]), .B(n41), .CO(n40), .S(sum[23]) );
  ADDHX1 U96 ( .A(a[18]), .B(n46), .CO(n45), .S(sum[18]) );
  ADDHX1 U97 ( .A(a[12]), .B(n52), .CO(n51), .S(sum[12]) );
  ADDHXL U98 ( .A(a[41]), .B(n23), .CO(n22), .S(sum[41]) );
  ADDHXL U99 ( .A(a[24]), .B(n40), .CO(n39), .S(sum[24]) );
  ADDHXL U100 ( .A(a[45]), .B(n19), .CO(n18), .S(sum[45]) );
  ADDHXL U101 ( .A(a[19]), .B(n45), .CO(n44), .S(sum[19]) );
  ADDHXL U102 ( .A(a[32]), .B(n32), .CO(n31), .S(sum[32]) );
  ADDHXL U103 ( .A(a[48]), .B(n16), .CO(n15), .S(sum[48]) );
  ADDHXL U104 ( .A(a[56]), .B(n8), .CO(n7), .S(sum[56]) );
  NOR2BX1 U105 ( .AN(a[60]), .B(n4), .Y(\sum[63] ) );
  ADDHXL U106 ( .A(a[49]), .B(n15), .CO(n14), .S(sum[49]) );
  ADDHXL U107 ( .A(a[11]), .B(n53), .CO(n52), .S(sum[11]) );
  ADDHXL U108 ( .A(a[17]), .B(n47), .CO(n46), .S(sum[17]) );
  ADDHXL U109 ( .A(a[30]), .B(n34), .CO(n33), .S(sum[30]) );
  ADDHXL U110 ( .A(a[38]), .B(n26), .CO(n25), .S(sum[38]) );
  ADDHXL U111 ( .A(a[22]), .B(n42), .CO(n41), .S(sum[22]) );
  ADDHXL U112 ( .A(a[28]), .B(n36), .CO(n35), .S(sum[28]) );
  ADDHXL U113 ( .A(a[2]), .B(n62), .CO(n61), .S(sum[2]) );
  ADDHXL U114 ( .A(a[10]), .B(n54), .CO(n53), .S(sum[10]) );
  ADDHXL U115 ( .A(a[20]), .B(n44), .CO(n43), .S(sum[20]) );
  ADDHXL U116 ( .A(a[8]), .B(n56), .CO(n55), .S(sum[8]) );
  ADDHXL U117 ( .A(a[59]), .B(n5), .CO(n4), .S(sum[59]) );
  ADDHXL U118 ( .A(a[4]), .B(n60), .CO(n59), .S(sum[4]) );
  ADDHXL U119 ( .A(a[33]), .B(n31), .CO(n30), .S(sum[33]) );
  ADDHXL U120 ( .A(a[43]), .B(n21), .CO(n20), .S(sum[43]) );
  ADDHXL U121 ( .A(a[51]), .B(n13), .CO(n12), .S(sum[51]) );
  ADDHXL U122 ( .A(a[13]), .B(n51), .CO(n50), .S(sum[13]) );
  ADDHXL U123 ( .A(a[57]), .B(n7), .CO(n6), .S(sum[57]) );
  ADDHXL U124 ( .A(carry_in), .B(a[0]), .CO(n63), .S(sum[0]) );
  XOR2X1 U125 ( .A(n4), .B(a[60]), .Y(sum[60]) );
endmodule


module GSIM_DW_div_tc_6 ( a, b, quotient, remainder, divide_by_0 );
  input [63:0] a;
  input [5:0] b;
  output [63:0] quotient;
  output [5:0] remainder;
  output divide_by_0;
  wire   \u_div/QInv[63] , \u_div/QInv[59] , \u_div/QInv[58] ,
         \u_div/QInv[57] , \u_div/QInv[56] , \u_div/QInv[55] ,
         \u_div/QInv[54] , \u_div/QInv[53] , \u_div/QInv[52] ,
         \u_div/QInv[51] , \u_div/QInv[50] , \u_div/QInv[49] ,
         \u_div/QInv[48] , \u_div/QInv[47] , \u_div/QInv[46] ,
         \u_div/QInv[45] , \u_div/QInv[44] , \u_div/QInv[43] ,
         \u_div/QInv[42] , \u_div/QInv[41] , \u_div/QInv[40] ,
         \u_div/QInv[39] , \u_div/QInv[38] , \u_div/QInv[37] ,
         \u_div/QInv[36] , \u_div/QInv[35] , \u_div/QInv[34] ,
         \u_div/QInv[33] , \u_div/QInv[32] , \u_div/QInv[31] ,
         \u_div/QInv[30] , \u_div/QInv[29] , \u_div/QInv[28] ,
         \u_div/QInv[27] , \u_div/QInv[26] , \u_div/QInv[25] ,
         \u_div/QInv[24] , \u_div/QInv[23] , \u_div/QInv[22] ,
         \u_div/QInv[21] , \u_div/QInv[20] , \u_div/QInv[19] ,
         \u_div/QInv[18] , \u_div/QInv[17] , \u_div/QInv[16] ,
         \u_div/QInv[15] , \u_div/QInv[14] , \u_div/QInv[13] ,
         \u_div/QInv[12] , \u_div/QInv[11] , \u_div/QInv[10] , \u_div/QInv[9] ,
         \u_div/QInv[8] , \u_div/QInv[7] , \u_div/QInv[6] , \u_div/QInv[5] ,
         \u_div/QInv[4] , \u_div/QInv[3] , \u_div/QInv[2] , \u_div/QInv[1] ,
         \u_div/QInv[0] , \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] ,
         \u_div/SumTmp[1][3] , \u_div/SumTmp[1][4] , \u_div/SumTmp[2][1] ,
         \u_div/SumTmp[2][2] , \u_div/SumTmp[2][3] , \u_div/SumTmp[2][4] ,
         \u_div/SumTmp[3][1] , \u_div/SumTmp[3][2] , \u_div/SumTmp[3][3] ,
         \u_div/SumTmp[3][4] , \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] ,
         \u_div/SumTmp[4][3] , \u_div/SumTmp[4][4] , \u_div/SumTmp[5][1] ,
         \u_div/SumTmp[5][2] , \u_div/SumTmp[5][3] , \u_div/SumTmp[5][4] ,
         \u_div/SumTmp[6][1] , \u_div/SumTmp[6][2] , \u_div/SumTmp[6][3] ,
         \u_div/SumTmp[6][4] , \u_div/SumTmp[7][1] , \u_div/SumTmp[7][2] ,
         \u_div/SumTmp[7][3] , \u_div/SumTmp[7][4] , \u_div/SumTmp[8][1] ,
         \u_div/SumTmp[8][2] , \u_div/SumTmp[8][3] , \u_div/SumTmp[8][4] ,
         \u_div/SumTmp[9][1] , \u_div/SumTmp[9][2] , \u_div/SumTmp[9][3] ,
         \u_div/SumTmp[9][4] , \u_div/SumTmp[10][1] , \u_div/SumTmp[10][2] ,
         \u_div/SumTmp[10][3] , \u_div/SumTmp[10][4] , \u_div/SumTmp[11][1] ,
         \u_div/SumTmp[11][2] , \u_div/SumTmp[11][3] , \u_div/SumTmp[11][4] ,
         \u_div/SumTmp[12][1] , \u_div/SumTmp[12][2] , \u_div/SumTmp[12][3] ,
         \u_div/SumTmp[12][4] , \u_div/SumTmp[13][1] , \u_div/SumTmp[13][2] ,
         \u_div/SumTmp[13][3] , \u_div/SumTmp[13][4] , \u_div/SumTmp[14][1] ,
         \u_div/SumTmp[14][2] , \u_div/SumTmp[14][3] , \u_div/SumTmp[14][4] ,
         \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] , \u_div/SumTmp[15][3] ,
         \u_div/SumTmp[15][4] , \u_div/SumTmp[16][1] , \u_div/SumTmp[16][2] ,
         \u_div/SumTmp[16][3] , \u_div/SumTmp[16][4] , \u_div/SumTmp[17][1] ,
         \u_div/SumTmp[17][2] , \u_div/SumTmp[17][3] , \u_div/SumTmp[17][4] ,
         \u_div/SumTmp[18][1] , \u_div/SumTmp[18][2] , \u_div/SumTmp[18][3] ,
         \u_div/SumTmp[18][4] , \u_div/SumTmp[19][1] , \u_div/SumTmp[19][2] ,
         \u_div/SumTmp[19][3] , \u_div/SumTmp[19][4] , \u_div/SumTmp[20][1] ,
         \u_div/SumTmp[20][2] , \u_div/SumTmp[20][3] , \u_div/SumTmp[20][4] ,
         \u_div/SumTmp[21][1] , \u_div/SumTmp[21][2] , \u_div/SumTmp[21][3] ,
         \u_div/SumTmp[21][4] , \u_div/SumTmp[22][1] , \u_div/SumTmp[22][2] ,
         \u_div/SumTmp[22][3] , \u_div/SumTmp[22][4] , \u_div/SumTmp[23][1] ,
         \u_div/SumTmp[23][2] , \u_div/SumTmp[23][3] , \u_div/SumTmp[23][4] ,
         \u_div/SumTmp[24][1] , \u_div/SumTmp[24][2] , \u_div/SumTmp[24][3] ,
         \u_div/SumTmp[24][4] , \u_div/SumTmp[25][1] , \u_div/SumTmp[25][2] ,
         \u_div/SumTmp[25][3] , \u_div/SumTmp[25][4] , \u_div/SumTmp[26][1] ,
         \u_div/SumTmp[26][2] , \u_div/SumTmp[26][3] , \u_div/SumTmp[26][4] ,
         \u_div/SumTmp[27][1] , \u_div/SumTmp[27][2] , \u_div/SumTmp[27][3] ,
         \u_div/SumTmp[27][4] , \u_div/SumTmp[28][1] , \u_div/SumTmp[28][2] ,
         \u_div/SumTmp[28][3] , \u_div/SumTmp[28][4] , \u_div/SumTmp[29][1] ,
         \u_div/SumTmp[29][2] , \u_div/SumTmp[29][3] , \u_div/SumTmp[29][4] ,
         \u_div/SumTmp[30][1] , \u_div/SumTmp[30][2] , \u_div/SumTmp[30][3] ,
         \u_div/SumTmp[30][4] , \u_div/SumTmp[31][1] , \u_div/SumTmp[31][2] ,
         \u_div/SumTmp[31][3] , \u_div/SumTmp[31][4] , \u_div/SumTmp[32][1] ,
         \u_div/SumTmp[32][2] , \u_div/SumTmp[32][3] , \u_div/SumTmp[32][4] ,
         \u_div/SumTmp[33][1] , \u_div/SumTmp[33][2] , \u_div/SumTmp[33][3] ,
         \u_div/SumTmp[33][4] , \u_div/SumTmp[34][1] , \u_div/SumTmp[34][2] ,
         \u_div/SumTmp[34][3] , \u_div/SumTmp[34][4] , \u_div/SumTmp[35][1] ,
         \u_div/SumTmp[35][2] , \u_div/SumTmp[35][3] , \u_div/SumTmp[35][4] ,
         \u_div/SumTmp[36][1] , \u_div/SumTmp[36][2] , \u_div/SumTmp[36][3] ,
         \u_div/SumTmp[36][4] , \u_div/SumTmp[37][1] , \u_div/SumTmp[37][2] ,
         \u_div/SumTmp[37][3] , \u_div/SumTmp[37][4] , \u_div/SumTmp[38][1] ,
         \u_div/SumTmp[38][2] , \u_div/SumTmp[38][3] , \u_div/SumTmp[38][4] ,
         \u_div/SumTmp[39][1] , \u_div/SumTmp[39][2] , \u_div/SumTmp[39][3] ,
         \u_div/SumTmp[39][4] , \u_div/SumTmp[40][1] , \u_div/SumTmp[40][2] ,
         \u_div/SumTmp[40][3] , \u_div/SumTmp[40][4] , \u_div/SumTmp[41][1] ,
         \u_div/SumTmp[41][2] , \u_div/SumTmp[41][3] , \u_div/SumTmp[41][4] ,
         \u_div/SumTmp[42][1] , \u_div/SumTmp[42][2] , \u_div/SumTmp[42][3] ,
         \u_div/SumTmp[42][4] , \u_div/SumTmp[43][1] , \u_div/SumTmp[43][2] ,
         \u_div/SumTmp[43][3] , \u_div/SumTmp[43][4] , \u_div/SumTmp[44][1] ,
         \u_div/SumTmp[44][2] , \u_div/SumTmp[44][3] , \u_div/SumTmp[44][4] ,
         \u_div/SumTmp[45][1] , \u_div/SumTmp[45][2] , \u_div/SumTmp[45][3] ,
         \u_div/SumTmp[45][4] , \u_div/SumTmp[46][1] , \u_div/SumTmp[46][2] ,
         \u_div/SumTmp[46][3] , \u_div/SumTmp[46][4] , \u_div/SumTmp[47][1] ,
         \u_div/SumTmp[47][2] , \u_div/SumTmp[47][3] , \u_div/SumTmp[47][4] ,
         \u_div/SumTmp[48][1] , \u_div/SumTmp[48][2] , \u_div/SumTmp[48][3] ,
         \u_div/SumTmp[48][4] , \u_div/SumTmp[49][1] , \u_div/SumTmp[49][2] ,
         \u_div/SumTmp[49][3] , \u_div/SumTmp[49][4] , \u_div/SumTmp[50][1] ,
         \u_div/SumTmp[50][2] , \u_div/SumTmp[50][3] , \u_div/SumTmp[50][4] ,
         \u_div/SumTmp[51][1] , \u_div/SumTmp[51][2] , \u_div/SumTmp[51][3] ,
         \u_div/SumTmp[51][4] , \u_div/SumTmp[52][1] , \u_div/SumTmp[52][2] ,
         \u_div/SumTmp[52][3] , \u_div/SumTmp[52][4] , \u_div/SumTmp[53][1] ,
         \u_div/SumTmp[53][2] , \u_div/SumTmp[53][3] , \u_div/SumTmp[53][4] ,
         \u_div/SumTmp[54][1] , \u_div/SumTmp[54][2] , \u_div/SumTmp[54][3] ,
         \u_div/SumTmp[54][4] , \u_div/SumTmp[55][1] , \u_div/SumTmp[55][2] ,
         \u_div/SumTmp[55][3] , \u_div/SumTmp[55][4] , \u_div/SumTmp[56][1] ,
         \u_div/SumTmp[56][2] , \u_div/SumTmp[56][3] , \u_div/SumTmp[56][4] ,
         \u_div/SumTmp[57][1] , \u_div/SumTmp[57][2] , \u_div/SumTmp[57][3] ,
         \u_div/SumTmp[57][4] , \u_div/SumTmp[58][1] , \u_div/SumTmp[58][2] ,
         \u_div/SumTmp[58][3] , \u_div/SumTmp[58][4] , \u_div/SumTmp[59][3] ,
         \u_div/SumTmp[59][4] , \u_div/CryTmp[0][6] , \u_div/CryTmp[1][6] ,
         \u_div/CryTmp[2][6] , \u_div/CryTmp[3][6] , \u_div/CryTmp[4][6] ,
         \u_div/CryTmp[5][6] , \u_div/CryTmp[6][6] , \u_div/CryTmp[7][6] ,
         \u_div/CryTmp[8][6] , \u_div/CryTmp[9][6] , \u_div/CryTmp[10][6] ,
         \u_div/CryTmp[11][6] , \u_div/CryTmp[12][6] , \u_div/CryTmp[13][6] ,
         \u_div/CryTmp[14][6] , \u_div/CryTmp[15][6] , \u_div/CryTmp[16][6] ,
         \u_div/CryTmp[17][6] , \u_div/CryTmp[18][6] , \u_div/CryTmp[19][6] ,
         \u_div/CryTmp[20][6] , \u_div/CryTmp[21][6] , \u_div/CryTmp[22][6] ,
         \u_div/CryTmp[23][6] , \u_div/CryTmp[24][6] , \u_div/CryTmp[25][6] ,
         \u_div/CryTmp[26][6] , \u_div/CryTmp[27][6] , \u_div/CryTmp[28][6] ,
         \u_div/CryTmp[29][6] , \u_div/CryTmp[30][6] , \u_div/CryTmp[31][6] ,
         \u_div/CryTmp[32][6] , \u_div/CryTmp[33][6] , \u_div/CryTmp[34][6] ,
         \u_div/CryTmp[35][6] , \u_div/CryTmp[36][6] , \u_div/CryTmp[37][6] ,
         \u_div/CryTmp[38][6] , \u_div/CryTmp[39][6] , \u_div/CryTmp[40][6] ,
         \u_div/CryTmp[41][6] , \u_div/CryTmp[42][6] , \u_div/CryTmp[43][6] ,
         \u_div/CryTmp[44][6] , \u_div/CryTmp[45][6] , \u_div/CryTmp[46][6] ,
         \u_div/CryTmp[47][6] , \u_div/CryTmp[48][6] , \u_div/CryTmp[49][6] ,
         \u_div/CryTmp[50][6] , \u_div/CryTmp[51][6] , \u_div/CryTmp[52][6] ,
         \u_div/CryTmp[53][6] , \u_div/CryTmp[54][6] , \u_div/CryTmp[55][6] ,
         \u_div/CryTmp[56][6] , \u_div/CryTmp[57][6] , \u_div/CryTmp[58][6] ,
         \u_div/CryTmp[59][6] , \u_div/PartRem[1][2] , \u_div/PartRem[1][3] ,
         \u_div/PartRem[1][4] , \u_div/PartRem[1][5] , \u_div/PartRem[2][2] ,
         \u_div/PartRem[2][3] , \u_div/PartRem[2][4] , \u_div/PartRem[2][5] ,
         \u_div/PartRem[3][0] , \u_div/PartRem[3][2] , \u_div/PartRem[3][3] ,
         \u_div/PartRem[3][4] , \u_div/PartRem[3][5] , \u_div/PartRem[4][0] ,
         \u_div/PartRem[4][2] , \u_div/PartRem[4][3] , \u_div/PartRem[4][4] ,
         \u_div/PartRem[4][5] , \u_div/PartRem[5][0] , \u_div/PartRem[5][2] ,
         \u_div/PartRem[5][3] , \u_div/PartRem[5][4] , \u_div/PartRem[5][5] ,
         \u_div/PartRem[6][0] , \u_div/PartRem[6][2] , \u_div/PartRem[6][3] ,
         \u_div/PartRem[6][4] , \u_div/PartRem[6][5] , \u_div/PartRem[7][0] ,
         \u_div/PartRem[7][2] , \u_div/PartRem[7][3] , \u_div/PartRem[7][4] ,
         \u_div/PartRem[7][5] , \u_div/PartRem[8][0] , \u_div/PartRem[8][2] ,
         \u_div/PartRem[8][3] , \u_div/PartRem[8][4] , \u_div/PartRem[8][5] ,
         \u_div/PartRem[9][0] , \u_div/PartRem[9][2] , \u_div/PartRem[9][3] ,
         \u_div/PartRem[9][4] , \u_div/PartRem[9][5] , \u_div/PartRem[10][0] ,
         \u_div/PartRem[10][2] , \u_div/PartRem[10][3] ,
         \u_div/PartRem[10][4] , \u_div/PartRem[10][5] ,
         \u_div/PartRem[11][0] , \u_div/PartRem[11][2] ,
         \u_div/PartRem[11][3] , \u_div/PartRem[11][4] ,
         \u_div/PartRem[11][5] , \u_div/PartRem[12][0] ,
         \u_div/PartRem[12][2] , \u_div/PartRem[12][3] ,
         \u_div/PartRem[12][4] , \u_div/PartRem[12][5] ,
         \u_div/PartRem[13][0] , \u_div/PartRem[13][2] ,
         \u_div/PartRem[13][3] , \u_div/PartRem[13][4] ,
         \u_div/PartRem[13][5] , \u_div/PartRem[14][0] ,
         \u_div/PartRem[14][2] , \u_div/PartRem[14][3] ,
         \u_div/PartRem[14][4] , \u_div/PartRem[14][5] ,
         \u_div/PartRem[15][0] , \u_div/PartRem[15][2] ,
         \u_div/PartRem[15][3] , \u_div/PartRem[15][4] ,
         \u_div/PartRem[15][5] , \u_div/PartRem[16][0] ,
         \u_div/PartRem[16][2] , \u_div/PartRem[16][3] ,
         \u_div/PartRem[16][4] , \u_div/PartRem[16][5] ,
         \u_div/PartRem[17][0] , \u_div/PartRem[17][2] ,
         \u_div/PartRem[17][3] , \u_div/PartRem[17][4] ,
         \u_div/PartRem[17][5] , \u_div/PartRem[18][0] ,
         \u_div/PartRem[18][2] , \u_div/PartRem[18][3] ,
         \u_div/PartRem[18][4] , \u_div/PartRem[18][5] ,
         \u_div/PartRem[19][0] , \u_div/PartRem[19][2] ,
         \u_div/PartRem[19][3] , \u_div/PartRem[19][4] ,
         \u_div/PartRem[19][5] , \u_div/PartRem[20][0] ,
         \u_div/PartRem[20][2] , \u_div/PartRem[20][3] ,
         \u_div/PartRem[20][4] , \u_div/PartRem[20][5] ,
         \u_div/PartRem[21][0] , \u_div/PartRem[21][2] ,
         \u_div/PartRem[21][3] , \u_div/PartRem[21][4] ,
         \u_div/PartRem[21][5] , \u_div/PartRem[22][0] ,
         \u_div/PartRem[22][2] , \u_div/PartRem[22][3] ,
         \u_div/PartRem[22][4] , \u_div/PartRem[22][5] ,
         \u_div/PartRem[23][0] , \u_div/PartRem[23][2] ,
         \u_div/PartRem[23][3] , \u_div/PartRem[23][4] ,
         \u_div/PartRem[23][5] , \u_div/PartRem[24][0] ,
         \u_div/PartRem[24][2] , \u_div/PartRem[24][3] ,
         \u_div/PartRem[24][4] , \u_div/PartRem[24][5] ,
         \u_div/PartRem[25][0] , \u_div/PartRem[25][2] ,
         \u_div/PartRem[25][3] , \u_div/PartRem[25][4] ,
         \u_div/PartRem[25][5] , \u_div/PartRem[26][0] ,
         \u_div/PartRem[26][2] , \u_div/PartRem[26][3] ,
         \u_div/PartRem[26][4] , \u_div/PartRem[26][5] ,
         \u_div/PartRem[27][0] , \u_div/PartRem[27][2] ,
         \u_div/PartRem[27][3] , \u_div/PartRem[27][4] ,
         \u_div/PartRem[27][5] , \u_div/PartRem[28][0] ,
         \u_div/PartRem[28][2] , \u_div/PartRem[28][3] ,
         \u_div/PartRem[28][4] , \u_div/PartRem[28][5] ,
         \u_div/PartRem[29][0] , \u_div/PartRem[29][2] ,
         \u_div/PartRem[29][3] , \u_div/PartRem[29][4] ,
         \u_div/PartRem[29][5] , \u_div/PartRem[30][0] ,
         \u_div/PartRem[30][2] , \u_div/PartRem[30][3] ,
         \u_div/PartRem[30][4] , \u_div/PartRem[30][5] ,
         \u_div/PartRem[31][0] , \u_div/PartRem[31][2] ,
         \u_div/PartRem[31][3] , \u_div/PartRem[31][4] ,
         \u_div/PartRem[31][5] , \u_div/PartRem[32][0] ,
         \u_div/PartRem[32][2] , \u_div/PartRem[32][3] ,
         \u_div/PartRem[32][4] , \u_div/PartRem[32][5] ,
         \u_div/PartRem[33][0] , \u_div/PartRem[33][2] ,
         \u_div/PartRem[33][3] , \u_div/PartRem[33][4] ,
         \u_div/PartRem[33][5] , \u_div/PartRem[34][0] ,
         \u_div/PartRem[34][2] , \u_div/PartRem[34][3] ,
         \u_div/PartRem[34][4] , \u_div/PartRem[34][5] ,
         \u_div/PartRem[35][0] , \u_div/PartRem[35][2] ,
         \u_div/PartRem[35][3] , \u_div/PartRem[35][4] ,
         \u_div/PartRem[35][5] , \u_div/PartRem[36][0] ,
         \u_div/PartRem[36][2] , \u_div/PartRem[36][3] ,
         \u_div/PartRem[36][4] , \u_div/PartRem[36][5] ,
         \u_div/PartRem[37][0] , \u_div/PartRem[37][2] ,
         \u_div/PartRem[37][3] , \u_div/PartRem[37][4] ,
         \u_div/PartRem[37][5] , \u_div/PartRem[38][0] ,
         \u_div/PartRem[38][2] , \u_div/PartRem[38][3] ,
         \u_div/PartRem[38][4] , \u_div/PartRem[38][5] ,
         \u_div/PartRem[39][0] , \u_div/PartRem[39][2] ,
         \u_div/PartRem[39][3] , \u_div/PartRem[39][4] ,
         \u_div/PartRem[39][5] , \u_div/PartRem[40][0] ,
         \u_div/PartRem[40][2] , \u_div/PartRem[40][3] ,
         \u_div/PartRem[40][4] , \u_div/PartRem[40][5] ,
         \u_div/PartRem[41][0] , \u_div/PartRem[41][2] ,
         \u_div/PartRem[41][3] , \u_div/PartRem[41][4] ,
         \u_div/PartRem[41][5] , \u_div/PartRem[42][0] ,
         \u_div/PartRem[42][2] , \u_div/PartRem[42][3] ,
         \u_div/PartRem[42][4] , \u_div/PartRem[42][5] ,
         \u_div/PartRem[43][0] , \u_div/PartRem[43][2] ,
         \u_div/PartRem[43][3] , \u_div/PartRem[43][4] ,
         \u_div/PartRem[43][5] , \u_div/PartRem[44][0] ,
         \u_div/PartRem[44][2] , \u_div/PartRem[44][3] ,
         \u_div/PartRem[44][4] , \u_div/PartRem[44][5] ,
         \u_div/PartRem[45][0] , \u_div/PartRem[45][2] ,
         \u_div/PartRem[45][3] , \u_div/PartRem[45][4] ,
         \u_div/PartRem[45][5] , \u_div/PartRem[46][0] ,
         \u_div/PartRem[46][2] , \u_div/PartRem[46][3] ,
         \u_div/PartRem[46][4] , \u_div/PartRem[46][5] ,
         \u_div/PartRem[47][0] , \u_div/PartRem[47][2] ,
         \u_div/PartRem[47][3] , \u_div/PartRem[47][4] ,
         \u_div/PartRem[47][5] , \u_div/PartRem[48][0] ,
         \u_div/PartRem[48][2] , \u_div/PartRem[48][3] ,
         \u_div/PartRem[48][4] , \u_div/PartRem[48][5] ,
         \u_div/PartRem[49][0] , \u_div/PartRem[49][2] ,
         \u_div/PartRem[49][3] , \u_div/PartRem[49][4] ,
         \u_div/PartRem[49][5] , \u_div/PartRem[50][0] ,
         \u_div/PartRem[50][2] , \u_div/PartRem[50][3] ,
         \u_div/PartRem[50][4] , \u_div/PartRem[50][5] ,
         \u_div/PartRem[51][0] , \u_div/PartRem[51][2] ,
         \u_div/PartRem[51][3] , \u_div/PartRem[51][4] ,
         \u_div/PartRem[51][5] , \u_div/PartRem[52][0] ,
         \u_div/PartRem[52][2] , \u_div/PartRem[52][3] ,
         \u_div/PartRem[52][4] , \u_div/PartRem[52][5] ,
         \u_div/PartRem[53][0] , \u_div/PartRem[53][2] ,
         \u_div/PartRem[53][3] , \u_div/PartRem[53][4] ,
         \u_div/PartRem[53][5] , \u_div/PartRem[54][0] ,
         \u_div/PartRem[54][2] , \u_div/PartRem[54][3] ,
         \u_div/PartRem[54][4] , \u_div/PartRem[54][5] ,
         \u_div/PartRem[55][0] , \u_div/PartRem[55][2] ,
         \u_div/PartRem[55][3] , \u_div/PartRem[55][4] ,
         \u_div/PartRem[55][5] , \u_div/PartRem[56][0] ,
         \u_div/PartRem[56][2] , \u_div/PartRem[56][3] ,
         \u_div/PartRem[56][4] , \u_div/PartRem[56][5] ,
         \u_div/PartRem[57][0] , \u_div/PartRem[57][2] ,
         \u_div/PartRem[57][3] , \u_div/PartRem[57][4] ,
         \u_div/PartRem[57][5] , \u_div/PartRem[58][0] ,
         \u_div/PartRem[58][2] , \u_div/PartRem[58][3] ,
         \u_div/PartRem[58][4] , \u_div/PartRem[58][5] ,
         \u_div/PartRem[59][0] , \u_div/PartRem[59][2] ,
         \u_div/PartRem[59][3] , \u_div/PartRem[59][4] ,
         \u_div/PartRem[59][5] , \u_div/PartRem[60][0] ,
         \u_div/PartRem[61][0] , \u_div/PartRem[62][0] ,
         \u_div/PartRem[63][0] , \u_div/PartRem[64][0] ,
         \u_div/u_add_PartRem_2_1/n3 , \u_div/u_add_PartRem_2_1/n2 ,
         \u_div/u_add_PartRem_2_2/n3 , \u_div/u_add_PartRem_2_2/n2 ,
         \u_div/u_add_PartRem_2_3/n3 , \u_div/u_add_PartRem_2_3/n2 ,
         \u_div/u_add_PartRem_2_4/n3 , \u_div/u_add_PartRem_2_4/n2 ,
         \u_div/u_add_PartRem_2_5/n3 , \u_div/u_add_PartRem_2_5/n2 ,
         \u_div/u_add_PartRem_2_6/n3 , \u_div/u_add_PartRem_2_6/n2 ,
         \u_div/u_add_PartRem_2_7/n3 , \u_div/u_add_PartRem_2_7/n2 ,
         \u_div/u_add_PartRem_2_8/n3 , \u_div/u_add_PartRem_2_8/n2 ,
         \u_div/u_add_PartRem_2_9/n3 , \u_div/u_add_PartRem_2_9/n2 ,
         \u_div/u_add_PartRem_2_10/n3 , \u_div/u_add_PartRem_2_10/n2 ,
         \u_div/u_add_PartRem_2_11/n3 , \u_div/u_add_PartRem_2_11/n2 ,
         \u_div/u_add_PartRem_2_12/n3 , \u_div/u_add_PartRem_2_12/n2 ,
         \u_div/u_add_PartRem_2_13/n3 , \u_div/u_add_PartRem_2_13/n2 ,
         \u_div/u_add_PartRem_2_14/n3 , \u_div/u_add_PartRem_2_14/n2 ,
         \u_div/u_add_PartRem_2_15/n3 , \u_div/u_add_PartRem_2_15/n2 ,
         \u_div/u_add_PartRem_2_16/n3 , \u_div/u_add_PartRem_2_16/n2 ,
         \u_div/u_add_PartRem_2_17/n3 , \u_div/u_add_PartRem_2_17/n2 ,
         \u_div/u_add_PartRem_2_18/n3 , \u_div/u_add_PartRem_2_18/n2 ,
         \u_div/u_add_PartRem_2_19/n3 , \u_div/u_add_PartRem_2_19/n2 ,
         \u_div/u_add_PartRem_2_20/n3 , \u_div/u_add_PartRem_2_20/n2 ,
         \u_div/u_add_PartRem_2_21/n3 , \u_div/u_add_PartRem_2_21/n2 ,
         \u_div/u_add_PartRem_2_22/n3 , \u_div/u_add_PartRem_2_22/n2 ,
         \u_div/u_add_PartRem_2_23/n3 , \u_div/u_add_PartRem_2_23/n2 ,
         \u_div/u_add_PartRem_2_24/n3 , \u_div/u_add_PartRem_2_24/n2 ,
         \u_div/u_add_PartRem_2_25/n3 , \u_div/u_add_PartRem_2_25/n2 ,
         \u_div/u_add_PartRem_2_26/n3 , \u_div/u_add_PartRem_2_26/n2 ,
         \u_div/u_add_PartRem_2_27/n3 , \u_div/u_add_PartRem_2_27/n2 ,
         \u_div/u_add_PartRem_2_28/n3 , \u_div/u_add_PartRem_2_28/n2 ,
         \u_div/u_add_PartRem_2_29/n3 , \u_div/u_add_PartRem_2_29/n2 ,
         \u_div/u_add_PartRem_2_30/n3 , \u_div/u_add_PartRem_2_30/n2 ,
         \u_div/u_add_PartRem_2_31/n3 , \u_div/u_add_PartRem_2_31/n2 ,
         \u_div/u_add_PartRem_2_32/n3 , \u_div/u_add_PartRem_2_32/n2 ,
         \u_div/u_add_PartRem_2_33/n3 , \u_div/u_add_PartRem_2_33/n2 ,
         \u_div/u_add_PartRem_2_34/n3 , \u_div/u_add_PartRem_2_34/n2 ,
         \u_div/u_add_PartRem_2_35/n3 , \u_div/u_add_PartRem_2_35/n2 ,
         \u_div/u_add_PartRem_2_36/n3 , \u_div/u_add_PartRem_2_36/n2 ,
         \u_div/u_add_PartRem_2_37/n3 , \u_div/u_add_PartRem_2_37/n2 ,
         \u_div/u_add_PartRem_2_38/n3 , \u_div/u_add_PartRem_2_38/n2 ,
         \u_div/u_add_PartRem_2_39/n3 , \u_div/u_add_PartRem_2_39/n2 ,
         \u_div/u_add_PartRem_2_40/n3 , \u_div/u_add_PartRem_2_40/n2 ,
         \u_div/u_add_PartRem_2_41/n3 , \u_div/u_add_PartRem_2_41/n2 ,
         \u_div/u_add_PartRem_2_42/n3 , \u_div/u_add_PartRem_2_42/n2 ,
         \u_div/u_add_PartRem_2_43/n3 , \u_div/u_add_PartRem_2_43/n2 ,
         \u_div/u_add_PartRem_2_44/n3 , \u_div/u_add_PartRem_2_44/n2 ,
         \u_div/u_add_PartRem_2_45/n3 , \u_div/u_add_PartRem_2_45/n2 ,
         \u_div/u_add_PartRem_2_46/n3 , \u_div/u_add_PartRem_2_46/n2 ,
         \u_div/u_add_PartRem_2_47/n3 , \u_div/u_add_PartRem_2_47/n2 ,
         \u_div/u_add_PartRem_2_48/n3 , \u_div/u_add_PartRem_2_48/n2 ,
         \u_div/u_add_PartRem_2_49/n3 , \u_div/u_add_PartRem_2_49/n2 ,
         \u_div/u_add_PartRem_2_50/n3 , \u_div/u_add_PartRem_2_50/n2 ,
         \u_div/u_add_PartRem_2_51/n3 , \u_div/u_add_PartRem_2_51/n2 ,
         \u_div/u_add_PartRem_2_52/n3 , \u_div/u_add_PartRem_2_52/n2 ,
         \u_div/u_add_PartRem_2_53/n3 , \u_div/u_add_PartRem_2_53/n2 ,
         \u_div/u_add_PartRem_2_54/n3 , \u_div/u_add_PartRem_2_54/n2 ,
         \u_div/u_add_PartRem_2_55/n3 , \u_div/u_add_PartRem_2_55/n2 ,
         \u_div/u_add_PartRem_2_56/n3 , \u_div/u_add_PartRem_2_56/n2 ,
         \u_div/u_add_PartRem_2_57/n3 , \u_div/u_add_PartRem_2_57/n2 ,
         \u_div/u_add_PartRem_2_58/n3 , \u_div/u_add_PartRem_2_58/n2 , n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign \u_div/QInv[63]  = a[63];

  GSIM_DW01_absval_6 \u_div/u_absval_AAbs  ( .A({n7, a[62:0]}), .ABSVAL({
        \u_div/PartRem[64][0] , \u_div/PartRem[63][0] , \u_div/PartRem[62][0] , 
        \u_div/PartRem[61][0] , \u_div/PartRem[60][0] , \u_div/PartRem[59][0] , 
        \u_div/PartRem[58][0] , \u_div/PartRem[57][0] , \u_div/PartRem[56][0] , 
        \u_div/PartRem[55][0] , \u_div/PartRem[54][0] , \u_div/PartRem[53][0] , 
        \u_div/PartRem[52][0] , \u_div/PartRem[51][0] , \u_div/PartRem[50][0] , 
        \u_div/PartRem[49][0] , \u_div/PartRem[48][0] , \u_div/PartRem[47][0] , 
        \u_div/PartRem[46][0] , \u_div/PartRem[45][0] , \u_div/PartRem[44][0] , 
        \u_div/PartRem[43][0] , \u_div/PartRem[42][0] , \u_div/PartRem[41][0] , 
        \u_div/PartRem[40][0] , \u_div/PartRem[39][0] , \u_div/PartRem[38][0] , 
        \u_div/PartRem[37][0] , \u_div/PartRem[36][0] , \u_div/PartRem[35][0] , 
        \u_div/PartRem[34][0] , \u_div/PartRem[33][0] , \u_div/PartRem[32][0] , 
        \u_div/PartRem[31][0] , \u_div/PartRem[30][0] , \u_div/PartRem[29][0] , 
        \u_div/PartRem[28][0] , \u_div/PartRem[27][0] , \u_div/PartRem[26][0] , 
        \u_div/PartRem[25][0] , \u_div/PartRem[24][0] , \u_div/PartRem[23][0] , 
        \u_div/PartRem[22][0] , \u_div/PartRem[21][0] , \u_div/PartRem[20][0] , 
        \u_div/PartRem[19][0] , \u_div/PartRem[18][0] , \u_div/PartRem[17][0] , 
        \u_div/PartRem[16][0] , \u_div/PartRem[15][0] , \u_div/PartRem[14][0] , 
        \u_div/PartRem[13][0] , \u_div/PartRem[12][0] , \u_div/PartRem[11][0] , 
        \u_div/PartRem[10][0] , \u_div/PartRem[9][0] , \u_div/PartRem[8][0] , 
        \u_div/PartRem[7][0] , \u_div/PartRem[6][0] , \u_div/PartRem[5][0] , 
        \u_div/PartRem[4][0] , \u_div/PartRem[3][0] , SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1}) );
  GSIM_DW_inc_6 \u_div/u_inc_QInc  ( .carry_in(n9), .a({n7, n7, n7, n8, 
        \u_div/QInv[59] , \u_div/QInv[58] , \u_div/QInv[57] , \u_div/QInv[56] , 
        \u_div/QInv[55] , \u_div/QInv[54] , \u_div/QInv[53] , \u_div/QInv[52] , 
        \u_div/QInv[51] , \u_div/QInv[50] , \u_div/QInv[49] , \u_div/QInv[48] , 
        \u_div/QInv[47] , \u_div/QInv[46] , \u_div/QInv[45] , \u_div/QInv[44] , 
        \u_div/QInv[43] , \u_div/QInv[42] , \u_div/QInv[41] , \u_div/QInv[40] , 
        \u_div/QInv[39] , \u_div/QInv[38] , \u_div/QInv[37] , \u_div/QInv[36] , 
        \u_div/QInv[35] , \u_div/QInv[34] , \u_div/QInv[33] , \u_div/QInv[32] , 
        \u_div/QInv[31] , \u_div/QInv[30] , \u_div/QInv[29] , \u_div/QInv[28] , 
        \u_div/QInv[27] , \u_div/QInv[26] , \u_div/QInv[25] , \u_div/QInv[24] , 
        \u_div/QInv[23] , \u_div/QInv[22] , \u_div/QInv[21] , \u_div/QInv[20] , 
        \u_div/QInv[19] , \u_div/QInv[18] , \u_div/QInv[17] , \u_div/QInv[16] , 
        \u_div/QInv[15] , \u_div/QInv[14] , \u_div/QInv[13] , \u_div/QInv[12] , 
        \u_div/QInv[11] , \u_div/QInv[10] , \u_div/QInv[9] , \u_div/QInv[8] , 
        \u_div/QInv[7] , \u_div/QInv[6] , \u_div/QInv[5] , \u_div/QInv[4] , 
        \u_div/QInv[3] , \u_div/QInv[2] , \u_div/QInv[1] , \u_div/QInv[0] }), 
        .sum(quotient) );
  ADDHXL \u_div/u_add_PartRem_2_7/U3  ( .A(\u_div/PartRem[8][4] ), .B(
        \u_div/u_add_PartRem_2_7/n3 ), .CO(\u_div/u_add_PartRem_2_7/n2 ), .S(
        \u_div/SumTmp[7][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_12/U3  ( .A(\u_div/PartRem[13][4] ), .B(
        \u_div/u_add_PartRem_2_12/n3 ), .CO(\u_div/u_add_PartRem_2_12/n2 ), 
        .S(\u_div/SumTmp[12][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_17/U3  ( .A(\u_div/PartRem[18][4] ), .B(
        \u_div/u_add_PartRem_2_17/n3 ), .CO(\u_div/u_add_PartRem_2_17/n2 ), 
        .S(\u_div/SumTmp[17][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_22/U3  ( .A(\u_div/PartRem[23][4] ), .B(
        \u_div/u_add_PartRem_2_22/n3 ), .CO(\u_div/u_add_PartRem_2_22/n2 ), 
        .S(\u_div/SumTmp[22][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_27/U3  ( .A(\u_div/PartRem[28][4] ), .B(
        \u_div/u_add_PartRem_2_27/n3 ), .CO(\u_div/u_add_PartRem_2_27/n2 ), 
        .S(\u_div/SumTmp[27][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_32/U3  ( .A(\u_div/PartRem[33][4] ), .B(
        \u_div/u_add_PartRem_2_32/n3 ), .CO(\u_div/u_add_PartRem_2_32/n2 ), 
        .S(\u_div/SumTmp[32][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_37/U3  ( .A(\u_div/PartRem[38][4] ), .B(
        \u_div/u_add_PartRem_2_37/n3 ), .CO(\u_div/u_add_PartRem_2_37/n2 ), 
        .S(\u_div/SumTmp[37][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_42/U3  ( .A(\u_div/PartRem[43][4] ), .B(
        \u_div/u_add_PartRem_2_42/n3 ), .CO(\u_div/u_add_PartRem_2_42/n2 ), 
        .S(\u_div/SumTmp[42][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_47/U3  ( .A(\u_div/PartRem[48][4] ), .B(
        \u_div/u_add_PartRem_2_47/n3 ), .CO(\u_div/u_add_PartRem_2_47/n2 ), 
        .S(\u_div/SumTmp[47][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_52/U3  ( .A(\u_div/PartRem[53][4] ), .B(
        \u_div/u_add_PartRem_2_52/n3 ), .CO(\u_div/u_add_PartRem_2_52/n2 ), 
        .S(\u_div/SumTmp[52][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_3_1  ( .A(\u_div/SumTmp[3][1] ), .B(
        \u_div/SumTmp[3][1] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_2_1  ( .A(\u_div/SumTmp[2][1] ), .B(
        \u_div/SumTmp[2][1] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_0  ( .A(\u_div/PartRem[7][0] ), .B(
        \u_div/PartRem[7][0] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/SumTmp[5][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_5_1  ( .A(\u_div/SumTmp[5][1] ), .B(
        \u_div/SumTmp[5][1] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_0  ( .A(\u_div/PartRem[12][0] ), .B(
        \u_div/PartRem[12][0] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/SumTmp[10][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_10_1  ( .A(\u_div/SumTmp[10][1] ), .B(
        \u_div/SumTmp[10][1] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_0  ( .A(\u_div/PartRem[17][0] ), .B(
        \u_div/PartRem[17][0] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/SumTmp[15][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_15_1  ( .A(\u_div/SumTmp[15][1] ), .B(
        \u_div/SumTmp[15][1] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_20_1  ( .A(\u_div/SumTmp[20][1] ), .B(
        \u_div/SumTmp[20][1] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_9_0  ( .A(\u_div/PartRem[10][0] ), .B(
        \u_div/PartRem[10][0] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/SumTmp[8][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_8_1  ( .A(\u_div/SumTmp[8][1] ), .B(
        \u_div/SumTmp[8][1] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_0  ( .A(\u_div/PartRem[15][0] ), .B(
        \u_div/PartRem[15][0] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/SumTmp[13][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_13_1  ( .A(\u_div/SumTmp[13][1] ), .B(
        \u_div/SumTmp[13][1] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_0  ( .A(\u_div/PartRem[20][0] ), .B(
        \u_div/PartRem[20][0] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/SumTmp[18][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_18_1  ( .A(\u_div/SumTmp[18][1] ), .B(
        \u_div/SumTmp[18][1] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_0  ( .A(\u_div/PartRem[25][0] ), .B(
        \u_div/PartRem[25][0] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/SumTmp[23][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_23_1  ( .A(\u_div/SumTmp[23][1] ), .B(
        \u_div/SumTmp[23][1] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_0  ( .A(\u_div/PartRem[8][0] ), .B(
        \u_div/PartRem[8][0] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/SumTmp[6][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_0  ( .A(\u_div/PartRem[13][0] ), .B(
        \u_div/PartRem[13][0] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/SumTmp[11][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_0  ( .A(\u_div/PartRem[18][0] ), .B(
        \u_div/PartRem[18][0] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/SumTmp[16][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_0  ( .A(\u_div/PartRem[23][0] ), .B(
        \u_div/PartRem[23][0] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/SumTmp[21][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_0  ( .A(\u_div/PartRem[26][0] ), .B(
        \u_div/PartRem[26][0] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/SumTmp[24][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_0  ( .A(\u_div/PartRem[27][0] ), .B(
        \u_div/PartRem[27][0] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/SumTmp[25][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_0  ( .A(\u_div/PartRem[28][0] ), .B(
        \u_div/PartRem[28][0] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/SumTmp[26][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_0  ( .A(\u_div/PartRem[29][0] ), .B(
        \u_div/PartRem[29][0] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/SumTmp[27][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_0  ( .A(\u_div/PartRem[31][0] ), .B(
        \u_div/PartRem[31][0] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/SumTmp[29][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_0  ( .A(\u_div/PartRem[32][0] ), .B(
        \u_div/PartRem[32][0] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/SumTmp[30][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_0  ( .A(\u_div/PartRem[33][0] ), .B(
        \u_div/PartRem[33][0] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/SumTmp[31][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_0  ( .A(\u_div/PartRem[34][0] ), .B(
        \u_div/PartRem[34][0] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/SumTmp[32][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_0  ( .A(\u_div/PartRem[36][0] ), .B(
        \u_div/PartRem[36][0] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/SumTmp[34][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_0  ( .A(\u_div/PartRem[37][0] ), .B(
        \u_div/PartRem[37][0] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/SumTmp[35][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_0  ( .A(\u_div/PartRem[38][0] ), .B(
        \u_div/PartRem[38][0] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/SumTmp[36][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_0  ( .A(\u_div/PartRem[39][0] ), .B(
        \u_div/PartRem[39][0] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/SumTmp[37][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_0  ( .A(\u_div/PartRem[41][0] ), .B(
        \u_div/PartRem[41][0] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/SumTmp[39][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_0  ( .A(\u_div/PartRem[42][0] ), .B(
        \u_div/PartRem[42][0] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/SumTmp[40][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_0  ( .A(\u_div/PartRem[43][0] ), .B(
        \u_div/PartRem[43][0] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/SumTmp[41][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_0  ( .A(\u_div/PartRem[44][0] ), .B(
        \u_div/PartRem[44][0] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/SumTmp[42][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_0  ( .A(\u_div/PartRem[46][0] ), .B(
        \u_div/PartRem[46][0] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/SumTmp[44][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_0  ( .A(\u_div/PartRem[47][0] ), .B(
        \u_div/PartRem[47][0] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/SumTmp[45][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_0  ( .A(\u_div/PartRem[48][0] ), .B(
        \u_div/PartRem[48][0] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/SumTmp[46][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_0  ( .A(\u_div/PartRem[49][0] ), .B(
        \u_div/PartRem[49][0] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/SumTmp[47][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_0  ( .A(\u_div/PartRem[51][0] ), .B(
        \u_div/PartRem[51][0] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/SumTmp[49][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_0  ( .A(\u_div/PartRem[52][0] ), .B(
        \u_div/PartRem[52][0] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/SumTmp[50][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_0  ( .A(\u_div/PartRem[53][0] ), .B(
        \u_div/PartRem[53][0] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/SumTmp[51][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_0  ( .A(\u_div/PartRem[54][0] ), .B(
        \u_div/PartRem[54][0] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/SumTmp[52][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_0  ( .A(\u_div/PartRem[56][0] ), .B(
        \u_div/PartRem[56][0] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/SumTmp[54][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_0  ( .A(\u_div/PartRem[57][0] ), .B(
        \u_div/PartRem[57][0] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/SumTmp[55][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_0  ( .A(\u_div/PartRem[58][0] ), .B(
        \u_div/PartRem[58][0] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/SumTmp[56][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_0  ( .A(\u_div/PartRem[59][0] ), .B(
        \u_div/PartRem[59][0] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/SumTmp[57][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_0  ( .A(\u_div/PartRem[60][0] ), .B(
        \u_div/PartRem[60][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/SumTmp[58][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_59_1  ( .A(\u_div/PartRem[61][0] ), .B(
        \u_div/PartRem[61][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_0  ( .A(\u_div/PartRem[30][0] ), .B(
        \u_div/PartRem[30][0] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/SumTmp[28][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_0  ( .A(\u_div/PartRem[35][0] ), .B(
        \u_div/PartRem[35][0] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/SumTmp[33][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_0  ( .A(\u_div/PartRem[40][0] ), .B(
        \u_div/PartRem[40][0] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/SumTmp[38][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_0  ( .A(\u_div/PartRem[45][0] ), .B(
        \u_div/PartRem[45][0] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/SumTmp[43][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_0  ( .A(\u_div/PartRem[50][0] ), .B(
        \u_div/PartRem[50][0] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/SumTmp[48][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_0  ( .A(\u_div/PartRem[55][0] ), .B(
        \u_div/PartRem[55][0] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/SumTmp[53][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_3  ( .A(\u_div/PartRem[29][3] ), .B(
        \u_div/SumTmp[28][3] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_3  ( .A(\u_div/PartRem[34][3] ), .B(
        \u_div/SumTmp[33][3] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_3  ( .A(\u_div/PartRem[39][3] ), .B(
        \u_div/SumTmp[38][3] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_3  ( .A(\u_div/PartRem[44][3] ), .B(
        \u_div/SumTmp[43][3] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_3  ( .A(\u_div/PartRem[49][3] ), .B(
        \u_div/SumTmp[48][3] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_3  ( .A(\u_div/PartRem[54][3] ), .B(
        \u_div/SumTmp[53][3] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_3  ( .A(\u_div/PartRem[8][3] ), .B(
        \u_div/SumTmp[7][3] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_3  ( .A(\u_div/PartRem[13][3] ), .B(
        \u_div/SumTmp[12][3] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_3  ( .A(\u_div/PartRem[18][3] ), .B(
        \u_div/SumTmp[17][3] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_3  ( .A(\u_div/PartRem[23][3] ), .B(
        \u_div/SumTmp[22][3] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_3  ( .A(\u_div/PartRem[26][3] ), .B(
        \u_div/SumTmp[25][3] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_3  ( .A(\u_div/PartRem[27][3] ), .B(
        \u_div/SumTmp[26][3] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_3  ( .A(\u_div/PartRem[28][3] ), .B(
        \u_div/SumTmp[27][3] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_3  ( .A(\u_div/PartRem[30][3] ), .B(
        \u_div/SumTmp[29][3] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_3  ( .A(\u_div/PartRem[31][3] ), .B(
        \u_div/SumTmp[30][3] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_3  ( .A(\u_div/PartRem[32][3] ), .B(
        \u_div/SumTmp[31][3] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_3  ( .A(\u_div/PartRem[33][3] ), .B(
        \u_div/SumTmp[32][3] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_3  ( .A(\u_div/PartRem[35][3] ), .B(
        \u_div/SumTmp[34][3] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_3  ( .A(\u_div/PartRem[36][3] ), .B(
        \u_div/SumTmp[35][3] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_3  ( .A(\u_div/PartRem[37][3] ), .B(
        \u_div/SumTmp[36][3] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_3  ( .A(\u_div/PartRem[38][3] ), .B(
        \u_div/SumTmp[37][3] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_3  ( .A(\u_div/PartRem[40][3] ), .B(
        \u_div/SumTmp[39][3] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_3  ( .A(\u_div/PartRem[41][3] ), .B(
        \u_div/SumTmp[40][3] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_3  ( .A(\u_div/PartRem[42][3] ), .B(
        \u_div/SumTmp[41][3] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_3  ( .A(\u_div/PartRem[43][3] ), .B(
        \u_div/SumTmp[42][3] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_3  ( .A(\u_div/PartRem[45][3] ), .B(
        \u_div/SumTmp[44][3] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_3  ( .A(\u_div/PartRem[46][3] ), .B(
        \u_div/SumTmp[45][3] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_3  ( .A(\u_div/PartRem[47][3] ), .B(
        \u_div/SumTmp[46][3] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_3  ( .A(\u_div/PartRem[48][3] ), .B(
        \u_div/SumTmp[47][3] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_3  ( .A(\u_div/PartRem[50][3] ), .B(
        \u_div/SumTmp[49][3] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_3  ( .A(\u_div/PartRem[51][3] ), .B(
        \u_div/SumTmp[50][3] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_3  ( .A(\u_div/PartRem[52][3] ), .B(
        \u_div/SumTmp[51][3] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_3  ( .A(\u_div/PartRem[53][3] ), .B(
        \u_div/SumTmp[52][3] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_3  ( .A(\u_div/PartRem[55][3] ), .B(
        \u_div/SumTmp[54][3] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_3  ( .A(\u_div/PartRem[56][3] ), .B(
        \u_div/SumTmp[55][3] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_3  ( .A(\u_div/PartRem[57][3] ), .B(
        \u_div/SumTmp[56][3] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_3  ( .A(\u_div/PartRem[58][3] ), .B(
        \u_div/SumTmp[57][3] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_3  ( .A(\u_div/PartRem[59][3] ), .B(
        \u_div/SumTmp[58][3] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_3  ( .A(\u_div/PartRem[63][0] ), .B(
        \u_div/SumTmp[59][3] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_1_1  ( .A(\u_div/SumTmp[1][1] ), .B(
        \u_div/SumTmp[1][1] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/SumTmp[1][2] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_2_4  ( .A(\u_div/PartRem[3][4] ), .B(
        \u_div/SumTmp[2][4] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_3_4  ( .A(\u_div/PartRem[4][4] ), .B(
        \u_div/SumTmp[3][4] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_9_4  ( .A(\u_div/PartRem[10][4] ), .B(
        \u_div/SumTmp[9][4] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_11_4  ( .A(\u_div/PartRem[12][4] ), .B(
        \u_div/SumTmp[11][4] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_21_4  ( .A(\u_div/PartRem[22][4] ), .B(
        \u_div/SumTmp[21][4] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_24_4  ( .A(\u_div/PartRem[25][4] ), .B(
        \u_div/SumTmp[24][4] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_5_4  ( .A(\u_div/PartRem[6][4] ), .B(
        \u_div/SumTmp[5][4] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_8_4  ( .A(\u_div/PartRem[9][4] ), .B(
        \u_div/SumTmp[8][4] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_10_4  ( .A(\u_div/PartRem[11][4] ), .B(
        \u_div/SumTmp[10][4] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_13_4  ( .A(\u_div/PartRem[14][4] ), .B(
        \u_div/SumTmp[13][4] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_15_4  ( .A(\u_div/PartRem[16][4] ), .B(
        \u_div/SumTmp[15][4] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_18_4  ( .A(\u_div/PartRem[19][4] ), .B(
        \u_div/SumTmp[18][4] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_20_4  ( .A(\u_div/PartRem[21][4] ), .B(
        \u_div/SumTmp[20][4] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_23_4  ( .A(\u_div/PartRem[24][4] ), .B(
        \u_div/SumTmp[23][4] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_4  ( .A(\u_div/PartRem[64][0] ), .B(
        \u_div/SumTmp[59][4] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_0  ( .A(\u_div/PartRem[3][0] ), .B(
        \u_div/PartRem[3][0] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/SumTmp[1][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_0  ( .A(\u_div/PartRem[4][0] ), .B(
        \u_div/PartRem[4][0] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/SumTmp[2][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_26_1  ( .A(\u_div/SumTmp[26][1] ), .B(
        \u_div/SumTmp[26][1] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_27_1  ( .A(\u_div/SumTmp[27][1] ), .B(
        \u_div/SumTmp[27][1] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_28_1  ( .A(\u_div/SumTmp[28][1] ), .B(
        \u_div/SumTmp[28][1] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_7_1  ( .A(\u_div/SumTmp[7][1] ), .B(
        \u_div/SumTmp[7][1] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_8_0  ( .A(\u_div/PartRem[9][0] ), .B(
        \u_div/PartRem[9][0] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/SumTmp[7][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_25_1  ( .A(\u_div/SumTmp[25][1] ), .B(
        \u_div/SumTmp[25][1] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_12_1  ( .A(\u_div/SumTmp[12][1] ), .B(
        \u_div/SumTmp[12][1] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_0  ( .A(\u_div/PartRem[14][0] ), .B(
        \u_div/PartRem[14][0] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/SumTmp[12][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_17_1  ( .A(\u_div/SumTmp[17][1] ), .B(
        \u_div/SumTmp[17][1] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_0  ( .A(\u_div/PartRem[19][0] ), .B(
        \u_div/PartRem[19][0] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/SumTmp[17][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_22_1  ( .A(\u_div/SumTmp[22][1] ), .B(
        \u_div/SumTmp[22][1] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_0  ( .A(\u_div/PartRem[24][0] ), .B(
        \u_div/PartRem[24][0] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/SumTmp[22][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_29_1  ( .A(\u_div/SumTmp[29][1] ), .B(
        \u_div/SumTmp[29][1] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_30_1  ( .A(\u_div/SumTmp[30][1] ), .B(
        \u_div/SumTmp[30][1] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_33_1  ( .A(\u_div/SumTmp[33][1] ), .B(
        \u_div/SumTmp[33][1] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_31_1  ( .A(\u_div/SumTmp[31][1] ), .B(
        \u_div/SumTmp[31][1] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_32_1  ( .A(\u_div/SumTmp[32][1] ), .B(
        \u_div/SumTmp[32][1] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_34_1  ( .A(\u_div/SumTmp[34][1] ), .B(
        \u_div/SumTmp[34][1] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_35_1  ( .A(\u_div/SumTmp[35][1] ), .B(
        \u_div/SumTmp[35][1] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_36_1  ( .A(\u_div/SumTmp[36][1] ), .B(
        \u_div/SumTmp[36][1] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_37_1  ( .A(\u_div/SumTmp[37][1] ), .B(
        \u_div/SumTmp[37][1] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_38_1  ( .A(\u_div/SumTmp[38][1] ), .B(
        \u_div/SumTmp[38][1] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_39_1  ( .A(\u_div/SumTmp[39][1] ), .B(
        \u_div/SumTmp[39][1] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_40_1  ( .A(\u_div/SumTmp[40][1] ), .B(
        \u_div/SumTmp[40][1] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_41_1  ( .A(\u_div/SumTmp[41][1] ), .B(
        \u_div/SumTmp[41][1] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_42_1  ( .A(\u_div/SumTmp[42][1] ), .B(
        \u_div/SumTmp[42][1] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_43_1  ( .A(\u_div/SumTmp[43][1] ), .B(
        \u_div/SumTmp[43][1] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_44_1  ( .A(\u_div/SumTmp[44][1] ), .B(
        \u_div/SumTmp[44][1] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_45_1  ( .A(\u_div/SumTmp[45][1] ), .B(
        \u_div/SumTmp[45][1] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_46_1  ( .A(\u_div/SumTmp[46][1] ), .B(
        \u_div/SumTmp[46][1] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_47_1  ( .A(\u_div/SumTmp[47][1] ), .B(
        \u_div/SumTmp[47][1] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_48_1  ( .A(\u_div/SumTmp[48][1] ), .B(
        \u_div/SumTmp[48][1] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_51_1  ( .A(\u_div/SumTmp[51][1] ), .B(
        \u_div/SumTmp[51][1] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_49_1  ( .A(\u_div/SumTmp[49][1] ), .B(
        \u_div/SumTmp[49][1] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_50_1  ( .A(\u_div/SumTmp[50][1] ), .B(
        \u_div/SumTmp[50][1] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_52_1  ( .A(\u_div/SumTmp[52][1] ), .B(
        \u_div/SumTmp[52][1] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_53_1  ( .A(\u_div/SumTmp[53][1] ), .B(
        \u_div/SumTmp[53][1] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_54_1  ( .A(\u_div/SumTmp[54][1] ), .B(
        \u_div/SumTmp[54][1] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_55_1  ( .A(\u_div/SumTmp[55][1] ), .B(
        \u_div/SumTmp[55][1] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_56_1  ( .A(\u_div/SumTmp[56][1] ), .B(
        \u_div/SumTmp[56][1] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_57_1  ( .A(\u_div/SumTmp[57][1] ), .B(
        \u_div/SumTmp[57][1] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_58_1  ( .A(\u_div/SumTmp[58][1] ), .B(
        \u_div/SumTmp[58][1] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_0  ( .A(\u_div/PartRem[6][0] ), .B(
        \u_div/PartRem[6][0] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/SumTmp[4][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_6_1  ( .A(\u_div/SumTmp[6][1] ), .B(
        \u_div/SumTmp[6][1] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_24_1  ( .A(\u_div/SumTmp[24][1] ), .B(
        \u_div/SumTmp[24][1] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_11_1  ( .A(\u_div/SumTmp[11][1] ), .B(
        \u_div/SumTmp[11][1] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_16_1  ( .A(\u_div/SumTmp[16][1] ), .B(
        \u_div/SumTmp[16][1] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_0  ( .A(\u_div/PartRem[11][0] ), .B(
        \u_div/PartRem[11][0] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/SumTmp[9][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_14_1  ( .A(\u_div/SumTmp[14][1] ), .B(
        \u_div/SumTmp[14][1] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_0  ( .A(\u_div/PartRem[16][0] ), .B(
        \u_div/PartRem[16][0] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/SumTmp[14][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_0  ( .A(\u_div/PartRem[21][0] ), .B(
        \u_div/PartRem[21][0] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/SumTmp[19][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_1_3  ( .A(\u_div/PartRem[2][3] ), .B(
        \u_div/SumTmp[1][3] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_2_3  ( .A(\u_div/PartRem[3][3] ), .B(
        \u_div/SumTmp[2][3] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_3_3  ( .A(\u_div/PartRem[4][3] ), .B(
        \u_div/SumTmp[3][3] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_5_3  ( .A(\u_div/PartRem[6][3] ), .B(
        \u_div/SumTmp[5][3] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_3  ( .A(\u_div/PartRem[11][3] ), .B(
        \u_div/SumTmp[10][3] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_15_3  ( .A(\u_div/PartRem[16][3] ), .B(
        \u_div/SumTmp[15][3] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_3  ( .A(\u_div/PartRem[21][3] ), .B(
        \u_div/SumTmp[20][3] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_8_3  ( .A(\u_div/PartRem[9][3] ), .B(
        \u_div/SumTmp[8][3] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_3  ( .A(\u_div/PartRem[14][3] ), .B(
        \u_div/SumTmp[13][3] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_3  ( .A(\u_div/PartRem[19][3] ), .B(
        \u_div/SumTmp[18][3] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_3  ( .A(\u_div/PartRem[24][3] ), .B(
        \u_div/SumTmp[23][3] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_3  ( .A(\u_div/PartRem[5][3] ), .B(
        \u_div/SumTmp[4][3] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_3  ( .A(\u_div/PartRem[7][3] ), .B(
        \u_div/SumTmp[6][3] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_3  ( .A(\u_div/PartRem[25][3] ), .B(
        \u_div/SumTmp[24][3] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_9_3  ( .A(\u_div/PartRem[10][3] ), .B(
        \u_div/SumTmp[9][3] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_3  ( .A(\u_div/PartRem[15][3] ), .B(
        \u_div/SumTmp[14][3] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_3  ( .A(\u_div/PartRem[20][3] ), .B(
        \u_div/SumTmp[19][3] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_11_3  ( .A(\u_div/PartRem[12][3] ), .B(
        \u_div/SumTmp[11][3] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_3  ( .A(\u_div/PartRem[17][3] ), .B(
        \u_div/SumTmp[16][3] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_3  ( .A(\u_div/PartRem[22][3] ), .B(
        \u_div/SumTmp[21][3] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_1_4  ( .A(\u_div/PartRem[2][4] ), .B(
        \u_div/SumTmp[1][4] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_4  ( .A(\u_div/PartRem[27][4] ), .B(
        \u_div/SumTmp[26][4] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_4  ( .A(\u_div/PartRem[29][4] ), .B(
        \u_div/SumTmp[28][4] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_4  ( .A(\u_div/PartRem[28][4] ), .B(
        \u_div/SumTmp[27][4] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_4  ( .A(\u_div/PartRem[34][4] ), .B(
        \u_div/SumTmp[33][4] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_4  ( .A(\u_div/PartRem[30][4] ), .B(
        \u_div/SumTmp[29][4] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_4  ( .A(\u_div/PartRem[31][4] ), .B(
        \u_div/SumTmp[30][4] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_4  ( .A(\u_div/PartRem[33][4] ), .B(
        \u_div/SumTmp[32][4] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_4  ( .A(\u_div/PartRem[32][4] ), .B(
        \u_div/SumTmp[31][4] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_4  ( .A(\u_div/PartRem[35][4] ), .B(
        \u_div/SumTmp[34][4] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_4  ( .A(\u_div/PartRem[39][4] ), .B(
        \u_div/SumTmp[38][4] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_4  ( .A(\u_div/PartRem[36][4] ), .B(
        \u_div/SumTmp[35][4] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_4  ( .A(\u_div/PartRem[37][4] ), .B(
        \u_div/SumTmp[36][4] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_4  ( .A(\u_div/PartRem[38][4] ), .B(
        \u_div/SumTmp[37][4] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_4  ( .A(\u_div/PartRem[40][4] ), .B(
        \u_div/SumTmp[39][4] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_4  ( .A(\u_div/PartRem[44][4] ), .B(
        \u_div/SumTmp[43][4] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_4  ( .A(\u_div/PartRem[41][4] ), .B(
        \u_div/SumTmp[40][4] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_4  ( .A(\u_div/PartRem[47][4] ), .B(
        \u_div/SumTmp[46][4] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_4  ( .A(\u_div/PartRem[42][4] ), .B(
        \u_div/SumTmp[41][4] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_4  ( .A(\u_div/PartRem[43][4] ), .B(
        \u_div/SumTmp[42][4] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_4  ( .A(\u_div/PartRem[50][4] ), .B(
        \u_div/SumTmp[49][4] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_4  ( .A(\u_div/PartRem[52][4] ), .B(
        \u_div/SumTmp[51][4] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_4  ( .A(\u_div/PartRem[46][4] ), .B(
        \u_div/SumTmp[45][4] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_4  ( .A(\u_div/PartRem[45][4] ), .B(
        \u_div/SumTmp[44][4] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_4  ( .A(\u_div/PartRem[49][4] ), .B(
        \u_div/SumTmp[48][4] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_4  ( .A(\u_div/PartRem[48][4] ), .B(
        \u_div/SumTmp[47][4] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_4  ( .A(\u_div/PartRem[51][4] ), .B(
        \u_div/SumTmp[50][4] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_4  ( .A(\u_div/PartRem[55][4] ), .B(
        \u_div/SumTmp[54][4] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_4  ( .A(\u_div/PartRem[53][4] ), .B(
        \u_div/SumTmp[52][4] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_4  ( .A(\u_div/PartRem[54][4] ), .B(
        \u_div/SumTmp[53][4] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_4  ( .A(\u_div/PartRem[58][4] ), .B(
        \u_div/SumTmp[57][4] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_4  ( .A(\u_div/PartRem[56][4] ), .B(
        \u_div/SumTmp[55][4] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_4  ( .A(\u_div/PartRem[57][4] ), .B(
        \u_div/SumTmp[56][4] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_4  ( .A(\u_div/PartRem[59][4] ), .B(
        \u_div/SumTmp[58][4] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_4  ( .A(\u_div/PartRem[8][4] ), .B(
        \u_div/SumTmp[7][4] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_4  ( .A(\u_div/PartRem[26][4] ), .B(
        \u_div/SumTmp[25][4] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_12_4  ( .A(\u_div/PartRem[13][4] ), .B(
        \u_div/SumTmp[12][4] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_4  ( .A(\u_div/PartRem[18][4] ), .B(
        \u_div/SumTmp[17][4] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_4  ( .A(\u_div/PartRem[23][4] ), .B(
        \u_div/SumTmp[22][4] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_14_4  ( .A(\u_div/PartRem[15][4] ), .B(
        \u_div/SumTmp[14][4] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][5] ) );
  MX2X6 \u_div/u_mx_PartRem_1_4_1  ( .A(\u_div/SumTmp[4][1] ), .B(
        \u_div/SumTmp[4][1] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][2] ) );
  CLKMX2X6 \u_div/u_mx_PartRem_1_9_1  ( .A(\u_div/SumTmp[9][1] ), .B(
        \u_div/SumTmp[9][1] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][2] ) );
  CLKMX2X6 \u_div/u_mx_PartRem_1_19_1  ( .A(\u_div/SumTmp[19][1] ), .B(
        \u_div/SumTmp[19][1] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_4  ( .A(\u_div/PartRem[20][4] ), .B(
        \u_div/SumTmp[19][4] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_6_4  ( .A(\u_div/PartRem[7][4] ), .B(
        \u_div/SumTmp[6][4] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_21_1  ( .A(\u_div/SumTmp[21][1] ), .B(
        \u_div/SumTmp[21][1] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][2] ) );
  MX2X1 \u_div/u_mx_PartRem_1_4_4  ( .A(\u_div/PartRem[5][4] ), .B(
        \u_div/SumTmp[4][4] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_0  ( .A(\u_div/PartRem[22][0] ), .B(
        \u_div/PartRem[22][0] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/SumTmp[20][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_0  ( .A(\u_div/PartRem[5][0] ), .B(
        \u_div/PartRem[5][0] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/SumTmp[3][1] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_4  ( .A(\u_div/PartRem[17][4] ), .B(
        \u_div/SumTmp[16][4] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][5] ) );
  OR2X6 U1 ( .A(\u_div/PartRem[17][5] ), .B(\u_div/u_add_PartRem_2_16/n2 ), 
        .Y(\u_div/CryTmp[16][6] ) );
  MXI2X2 U2 ( .A(\u_div/SumTmp[21][2] ), .B(\u_div/PartRem[22][2] ), .S0(
        \u_div/CryTmp[21][6] ), .Y(\u_div/PartRem[21][3] ) );
  ADDHXL U3 ( .A(\u_div/PartRem[14][4] ), .B(\u_div/u_add_PartRem_2_13/n3 ), 
        .CO(\u_div/u_add_PartRem_2_13/n2 ), .S(\u_div/SumTmp[13][4] ) );
  ADDHXL U4 ( .A(\u_div/PartRem[19][4] ), .B(\u_div/u_add_PartRem_2_18/n3 ), 
        .CO(\u_div/u_add_PartRem_2_18/n2 ), .S(\u_div/SumTmp[18][4] ) );
  ADDHXL U5 ( .A(\u_div/PartRem[9][4] ), .B(\u_div/u_add_PartRem_2_8/n3 ), 
        .CO(\u_div/u_add_PartRem_2_8/n2 ), .S(\u_div/SumTmp[8][4] ) );
  NOR2X1 U6 ( .A(\u_div/PartRem[63][0] ), .B(\u_div/PartRem[62][0] ), .Y(n12)
         );
  OR2X6 U7 ( .A(\u_div/PartRem[20][5] ), .B(\u_div/u_add_PartRem_2_19/n2 ), 
        .Y(\u_div/CryTmp[19][6] ) );
  OR2X6 U8 ( .A(\u_div/PartRem[10][5] ), .B(\u_div/u_add_PartRem_2_9/n2 ), .Y(
        \u_div/CryTmp[9][6] ) );
  OR2X6 U9 ( .A(\u_div/PartRem[5][5] ), .B(\u_div/u_add_PartRem_2_4/n2 ), .Y(
        \u_div/CryTmp[4][6] ) );
  OR2X2 U10 ( .A(\u_div/PartRem[7][5] ), .B(\u_div/u_add_PartRem_2_6/n2 ), .Y(
        \u_div/CryTmp[6][6] ) );
  XOR2XL U11 ( .A(\u_div/CryTmp[19][6] ), .B(n7), .Y(\u_div/QInv[19] ) );
  MXI2X4 U12 ( .A(\u_div/SumTmp[19][2] ), .B(\u_div/PartRem[20][2] ), .S0(
        \u_div/CryTmp[19][6] ), .Y(\u_div/PartRem[19][3] ) );
  XOR2XL U13 ( .A(\u_div/CryTmp[9][6] ), .B(n7), .Y(\u_div/QInv[9] ) );
  MXI2X4 U14 ( .A(\u_div/SumTmp[9][2] ), .B(\u_div/PartRem[10][2] ), .S0(
        \u_div/CryTmp[9][6] ), .Y(\u_div/PartRem[9][3] ) );
  XOR2XL U15 ( .A(\u_div/CryTmp[4][6] ), .B(n9), .Y(\u_div/QInv[4] ) );
  MXI2X4 U16 ( .A(\u_div/SumTmp[4][2] ), .B(\u_div/PartRem[5][2] ), .S0(
        \u_div/CryTmp[4][6] ), .Y(\u_div/PartRem[4][3] ) );
  XOR2XL U17 ( .A(\u_div/CryTmp[21][6] ), .B(n7), .Y(\u_div/QInv[21] ) );
  OR2X6 U18 ( .A(\u_div/PartRem[22][5] ), .B(\u_div/u_add_PartRem_2_21/n2 ), 
        .Y(\u_div/CryTmp[21][6] ) );
  OR2X8 U19 ( .A(\u_div/PartRem[12][5] ), .B(\u_div/u_add_PartRem_2_11/n2 ), 
        .Y(\u_div/CryTmp[11][6] ) );
  ADDHX2 U20 ( .A(\u_div/PartRem[12][4] ), .B(\u_div/u_add_PartRem_2_11/n3 ), 
        .CO(\u_div/u_add_PartRem_2_11/n2 ), .S(\u_div/SumTmp[11][4] ) );
  OR2X6 U21 ( .A(\u_div/PartRem[4][5] ), .B(\u_div/u_add_PartRem_2_3/n2 ), .Y(
        \u_div/CryTmp[3][6] ) );
  OR2X1 U22 ( .A(\u_div/PartRem[14][5] ), .B(\u_div/u_add_PartRem_2_13/n2 ), 
        .Y(\u_div/CryTmp[13][6] ) );
  OR2X1 U23 ( .A(\u_div/PartRem[19][5] ), .B(\u_div/u_add_PartRem_2_18/n2 ), 
        .Y(\u_div/CryTmp[18][6] ) );
  OR2X1 U24 ( .A(\u_div/PartRem[9][5] ), .B(\u_div/u_add_PartRem_2_8/n2 ), .Y(
        \u_div/CryTmp[8][6] ) );
  ADDHXL U25 ( .A(\u_div/PartRem[58][4] ), .B(\u_div/u_add_PartRem_2_57/n3 ), 
        .CO(\u_div/u_add_PartRem_2_57/n2 ), .S(\u_div/SumTmp[57][4] ) );
  ADDHXL U26 ( .A(\u_div/PartRem[57][4] ), .B(\u_div/u_add_PartRem_2_56/n3 ), 
        .CO(\u_div/u_add_PartRem_2_56/n2 ), .S(\u_div/SumTmp[56][4] ) );
  ADDHXL U27 ( .A(\u_div/PartRem[56][4] ), .B(\u_div/u_add_PartRem_2_55/n3 ), 
        .CO(\u_div/u_add_PartRem_2_55/n2 ), .S(\u_div/SumTmp[55][4] ) );
  ADDHXL U28 ( .A(\u_div/PartRem[55][4] ), .B(\u_div/u_add_PartRem_2_54/n3 ), 
        .CO(\u_div/u_add_PartRem_2_54/n2 ), .S(\u_div/SumTmp[54][4] ) );
  ADDHXL U29 ( .A(\u_div/PartRem[51][4] ), .B(\u_div/u_add_PartRem_2_50/n3 ), 
        .CO(\u_div/u_add_PartRem_2_50/n2 ), .S(\u_div/SumTmp[50][4] ) );
  ADDHXL U30 ( .A(\u_div/PartRem[50][4] ), .B(\u_div/u_add_PartRem_2_49/n3 ), 
        .CO(\u_div/u_add_PartRem_2_49/n2 ), .S(\u_div/SumTmp[49][4] ) );
  ADDHXL U31 ( .A(\u_div/PartRem[49][4] ), .B(\u_div/u_add_PartRem_2_48/n3 ), 
        .CO(\u_div/u_add_PartRem_2_48/n2 ), .S(\u_div/SumTmp[48][4] ) );
  ADDHXL U32 ( .A(\u_div/PartRem[47][4] ), .B(\u_div/u_add_PartRem_2_46/n3 ), 
        .CO(\u_div/u_add_PartRem_2_46/n2 ), .S(\u_div/SumTmp[46][4] ) );
  ADDHXL U33 ( .A(\u_div/PartRem[42][4] ), .B(\u_div/u_add_PartRem_2_41/n3 ), 
        .CO(\u_div/u_add_PartRem_2_41/n2 ), .S(\u_div/SumTmp[41][4] ) );
  ADDHXL U34 ( .A(\u_div/PartRem[41][4] ), .B(\u_div/u_add_PartRem_2_40/n3 ), 
        .CO(\u_div/u_add_PartRem_2_40/n2 ), .S(\u_div/SumTmp[40][4] ) );
  ADDHXL U35 ( .A(\u_div/PartRem[40][4] ), .B(\u_div/u_add_PartRem_2_39/n3 ), 
        .CO(\u_div/u_add_PartRem_2_39/n2 ), .S(\u_div/SumTmp[39][4] ) );
  ADDHXL U36 ( .A(\u_div/PartRem[39][4] ), .B(\u_div/u_add_PartRem_2_38/n3 ), 
        .CO(\u_div/u_add_PartRem_2_38/n2 ), .S(\u_div/SumTmp[38][4] ) );
  ADDHXL U37 ( .A(\u_div/PartRem[37][4] ), .B(\u_div/u_add_PartRem_2_36/n3 ), 
        .CO(\u_div/u_add_PartRem_2_36/n2 ), .S(\u_div/SumTmp[36][4] ) );
  ADDHXL U38 ( .A(\u_div/PartRem[32][4] ), .B(\u_div/u_add_PartRem_2_31/n3 ), 
        .CO(\u_div/u_add_PartRem_2_31/n2 ), .S(\u_div/SumTmp[31][4] ) );
  ADDHXL U39 ( .A(\u_div/PartRem[31][4] ), .B(\u_div/u_add_PartRem_2_30/n3 ), 
        .CO(\u_div/u_add_PartRem_2_30/n2 ), .S(\u_div/SumTmp[30][4] ) );
  ADDHXL U40 ( .A(\u_div/PartRem[30][4] ), .B(\u_div/u_add_PartRem_2_29/n3 ), 
        .CO(\u_div/u_add_PartRem_2_29/n2 ), .S(\u_div/SumTmp[29][4] ) );
  ADDHXL U41 ( .A(\u_div/PartRem[29][4] ), .B(\u_div/u_add_PartRem_2_28/n3 ), 
        .CO(\u_div/u_add_PartRem_2_28/n2 ), .S(\u_div/SumTmp[28][4] ) );
  ADDHXL U42 ( .A(\u_div/PartRem[27][4] ), .B(\u_div/u_add_PartRem_2_26/n3 ), 
        .CO(\u_div/u_add_PartRem_2_26/n2 ), .S(\u_div/SumTmp[26][4] ) );
  ADDHXL U43 ( .A(\u_div/PartRem[54][4] ), .B(\u_div/u_add_PartRem_2_53/n3 ), 
        .CO(\u_div/u_add_PartRem_2_53/n2 ), .S(\u_div/SumTmp[53][4] ) );
  ADDHXL U44 ( .A(\u_div/PartRem[52][4] ), .B(\u_div/u_add_PartRem_2_51/n3 ), 
        .CO(\u_div/u_add_PartRem_2_51/n2 ), .S(\u_div/SumTmp[51][4] ) );
  ADDHXL U45 ( .A(\u_div/PartRem[46][4] ), .B(\u_div/u_add_PartRem_2_45/n3 ), 
        .CO(\u_div/u_add_PartRem_2_45/n2 ), .S(\u_div/SumTmp[45][4] ) );
  ADDHXL U46 ( .A(\u_div/PartRem[45][4] ), .B(\u_div/u_add_PartRem_2_44/n3 ), 
        .CO(\u_div/u_add_PartRem_2_44/n2 ), .S(\u_div/SumTmp[44][4] ) );
  ADDHXL U47 ( .A(\u_div/PartRem[44][4] ), .B(\u_div/u_add_PartRem_2_43/n3 ), 
        .CO(\u_div/u_add_PartRem_2_43/n2 ), .S(\u_div/SumTmp[43][4] ) );
  ADDHXL U48 ( .A(\u_div/PartRem[36][4] ), .B(\u_div/u_add_PartRem_2_35/n3 ), 
        .CO(\u_div/u_add_PartRem_2_35/n2 ), .S(\u_div/SumTmp[35][4] ) );
  ADDHXL U49 ( .A(\u_div/PartRem[35][4] ), .B(\u_div/u_add_PartRem_2_34/n3 ), 
        .CO(\u_div/u_add_PartRem_2_34/n2 ), .S(\u_div/SumTmp[34][4] ) );
  ADDHXL U50 ( .A(\u_div/PartRem[34][4] ), .B(\u_div/u_add_PartRem_2_33/n3 ), 
        .CO(\u_div/u_add_PartRem_2_33/n2 ), .S(\u_div/SumTmp[33][4] ) );
  ADDHXL U51 ( .A(\u_div/PartRem[26][4] ), .B(\u_div/u_add_PartRem_2_25/n3 ), 
        .CO(\u_div/u_add_PartRem_2_25/n2 ), .S(\u_div/SumTmp[25][4] ) );
  ADDHXL U52 ( .A(\u_div/PartRem[25][4] ), .B(\u_div/u_add_PartRem_2_24/n3 ), 
        .CO(\u_div/u_add_PartRem_2_24/n2 ), .S(\u_div/SumTmp[24][4] ) );
  ADDHXL U53 ( .A(\u_div/PartRem[22][4] ), .B(\u_div/u_add_PartRem_2_21/n3 ), 
        .CO(\u_div/u_add_PartRem_2_21/n2 ), .S(\u_div/SumTmp[21][4] ) );
  ADDHXL U54 ( .A(\u_div/PartRem[17][4] ), .B(\u_div/u_add_PartRem_2_16/n3 ), 
        .CO(\u_div/u_add_PartRem_2_16/n2 ), .S(\u_div/SumTmp[16][4] ) );
  ADDHXL U55 ( .A(\u_div/PartRem[7][4] ), .B(\u_div/u_add_PartRem_2_6/n3 ), 
        .CO(\u_div/u_add_PartRem_2_6/n2 ), .S(\u_div/SumTmp[6][4] ) );
  ADDHXL U56 ( .A(\u_div/PartRem[15][4] ), .B(\u_div/u_add_PartRem_2_14/n3 ), 
        .CO(\u_div/u_add_PartRem_2_14/n2 ), .S(\u_div/SumTmp[14][4] ) );
  INVXL U57 ( .A(\u_div/PartRem[20][2] ), .Y(\u_div/SumTmp[19][2] ) );
  INVXL U58 ( .A(\u_div/PartRem[10][2] ), .Y(\u_div/SumTmp[9][2] ) );
  INVXL U59 ( .A(\u_div/PartRem[5][2] ), .Y(\u_div/SumTmp[4][2] ) );
  INVXL U60 ( .A(\u_div/PartRem[15][2] ), .Y(\u_div/SumTmp[14][2] ) );
  INVXL U61 ( .A(\u_div/PartRem[3][2] ), .Y(\u_div/SumTmp[2][2] ) );
  NOR2BX4 U62 ( .AN(\u_div/PartRem[64][0] ), .B(n12), .Y(\u_div/CryTmp[59][6] ) );
  NAND2BX4 U63 ( .AN(\u_div/PartRem[11][5] ), .B(n3), .Y(\u_div/CryTmp[10][6] ) );
  INVX3 U64 ( .A(\u_div/u_add_PartRem_2_10/n2 ), .Y(n3) );
  NAND2BX4 U65 ( .AN(\u_div/PartRem[16][5] ), .B(n2), .Y(\u_div/CryTmp[15][6] ) );
  INVX3 U66 ( .A(\u_div/u_add_PartRem_2_15/n2 ), .Y(n2) );
  NAND2BX4 U67 ( .AN(\u_div/PartRem[21][5] ), .B(n1), .Y(\u_div/CryTmp[20][6] ) );
  INVX3 U68 ( .A(\u_div/u_add_PartRem_2_20/n2 ), .Y(n1) );
  NAND2BX4 U69 ( .AN(\u_div/PartRem[6][5] ), .B(n5), .Y(\u_div/CryTmp[5][6] )
         );
  INVX3 U70 ( .A(\u_div/u_add_PartRem_2_5/n2 ), .Y(n5) );
  NAND2BX4 U71 ( .AN(\u_div/PartRem[24][5] ), .B(n4), .Y(\u_div/CryTmp[23][6] ) );
  INVX3 U72 ( .A(\u_div/u_add_PartRem_2_23/n2 ), .Y(n4) );
  MXI2X2 U73 ( .A(\u_div/SumTmp[11][2] ), .B(\u_div/PartRem[12][2] ), .S0(
        \u_div/CryTmp[11][6] ), .Y(\u_div/PartRem[11][3] ) );
  MXI2X2 U74 ( .A(\u_div/SumTmp[24][2] ), .B(\u_div/PartRem[25][2] ), .S0(
        \u_div/CryTmp[24][6] ), .Y(\u_div/PartRem[24][3] ) );
  MXI2X2 U75 ( .A(\u_div/SumTmp[14][2] ), .B(\u_div/PartRem[15][2] ), .S0(
        \u_div/CryTmp[14][6] ), .Y(\u_div/PartRem[14][3] ) );
  MXI2X2 U76 ( .A(\u_div/SumTmp[16][2] ), .B(\u_div/PartRem[17][2] ), .S0(
        \u_div/CryTmp[16][6] ), .Y(\u_div/PartRem[16][3] ) );
  MXI2X2 U77 ( .A(\u_div/SumTmp[6][2] ), .B(\u_div/PartRem[7][2] ), .S0(
        \u_div/CryTmp[6][6] ), .Y(\u_div/PartRem[6][3] ) );
  MXI2X2 U78 ( .A(\u_div/SumTmp[28][2] ), .B(\u_div/PartRem[29][2] ), .S0(
        \u_div/CryTmp[28][6] ), .Y(\u_div/PartRem[28][3] ) );
  MXI2X2 U79 ( .A(\u_div/SumTmp[2][2] ), .B(\u_div/PartRem[3][2] ), .S0(
        \u_div/CryTmp[2][6] ), .Y(\u_div/PartRem[2][3] ) );
  ADDHX1 U80 ( .A(\u_div/PartRem[3][4] ), .B(\u_div/u_add_PartRem_2_2/n3 ), 
        .CO(\u_div/u_add_PartRem_2_2/n2 ), .S(\u_div/SumTmp[2][4] ) );
  OR2X2 U81 ( .A(\u_div/PartRem[3][2] ), .B(\u_div/PartRem[3][3] ), .Y(
        \u_div/u_add_PartRem_2_2/n3 ) );
  ADDHX1 U82 ( .A(\u_div/PartRem[5][4] ), .B(\u_div/u_add_PartRem_2_4/n3 ), 
        .CO(\u_div/u_add_PartRem_2_4/n2 ), .S(\u_div/SumTmp[4][4] ) );
  OR2X2 U83 ( .A(\u_div/PartRem[5][2] ), .B(\u_div/PartRem[5][3] ), .Y(
        \u_div/u_add_PartRem_2_4/n3 ) );
  OR2X2 U84 ( .A(\u_div/PartRem[17][2] ), .B(\u_div/PartRem[17][3] ), .Y(
        \u_div/u_add_PartRem_2_16/n3 ) );
  OR2X2 U85 ( .A(\u_div/PartRem[22][2] ), .B(\u_div/PartRem[22][3] ), .Y(
        \u_div/u_add_PartRem_2_21/n3 ) );
  OR2X2 U86 ( .A(\u_div/PartRem[7][2] ), .B(\u_div/PartRem[7][3] ), .Y(
        \u_div/u_add_PartRem_2_6/n3 ) );
  OR2X2 U87 ( .A(\u_div/PartRem[12][2] ), .B(\u_div/PartRem[12][3] ), .Y(
        \u_div/u_add_PartRem_2_11/n3 ) );
  OR2X2 U88 ( .A(\u_div/PartRem[25][2] ), .B(\u_div/PartRem[25][3] ), .Y(
        \u_div/u_add_PartRem_2_24/n3 ) );
  ADDHX1 U89 ( .A(\u_div/PartRem[10][4] ), .B(\u_div/u_add_PartRem_2_9/n3 ), 
        .CO(\u_div/u_add_PartRem_2_9/n2 ), .S(\u_div/SumTmp[9][4] ) );
  OR2X2 U90 ( .A(\u_div/PartRem[10][2] ), .B(\u_div/PartRem[10][3] ), .Y(
        \u_div/u_add_PartRem_2_9/n3 ) );
  ADDHX1 U91 ( .A(\u_div/PartRem[20][4] ), .B(\u_div/u_add_PartRem_2_19/n3 ), 
        .CO(\u_div/u_add_PartRem_2_19/n2 ), .S(\u_div/SumTmp[19][4] ) );
  OR2X2 U92 ( .A(\u_div/PartRem[20][2] ), .B(\u_div/PartRem[20][3] ), .Y(
        \u_div/u_add_PartRem_2_19/n3 ) );
  OR2X2 U93 ( .A(\u_div/PartRem[26][2] ), .B(\u_div/PartRem[26][3] ), .Y(
        \u_div/u_add_PartRem_2_25/n3 ) );
  OR2X2 U94 ( .A(\u_div/PartRem[27][2] ), .B(\u_div/PartRem[27][3] ), .Y(
        \u_div/u_add_PartRem_2_26/n3 ) );
  OR2X2 U95 ( .A(\u_div/PartRem[29][2] ), .B(\u_div/PartRem[29][3] ), .Y(
        \u_div/u_add_PartRem_2_28/n3 ) );
  OR2X2 U96 ( .A(\u_div/PartRem[34][2] ), .B(\u_div/PartRem[34][3] ), .Y(
        \u_div/u_add_PartRem_2_33/n3 ) );
  OR2X2 U97 ( .A(\u_div/PartRem[42][2] ), .B(\u_div/PartRem[42][3] ), .Y(
        \u_div/u_add_PartRem_2_41/n3 ) );
  OR2X2 U98 ( .A(\u_div/PartRem[35][2] ), .B(\u_div/PartRem[35][3] ), .Y(
        \u_div/u_add_PartRem_2_34/n3 ) );
  OR2X2 U99 ( .A(\u_div/PartRem[39][2] ), .B(\u_div/PartRem[39][3] ), .Y(
        \u_div/u_add_PartRem_2_38/n3 ) );
  OR2X2 U100 ( .A(\u_div/PartRem[41][2] ), .B(\u_div/PartRem[41][3] ), .Y(
        \u_div/u_add_PartRem_2_40/n3 ) );
  OR2X2 U101 ( .A(\u_div/PartRem[36][2] ), .B(\u_div/PartRem[36][3] ), .Y(
        \u_div/u_add_PartRem_2_35/n3 ) );
  OR2X2 U102 ( .A(\u_div/PartRem[30][2] ), .B(\u_div/PartRem[30][3] ), .Y(
        \u_div/u_add_PartRem_2_29/n3 ) );
  OR2X2 U103 ( .A(\u_div/PartRem[32][2] ), .B(\u_div/PartRem[32][3] ), .Y(
        \u_div/u_add_PartRem_2_31/n3 ) );
  OR2X2 U104 ( .A(\u_div/PartRem[44][2] ), .B(\u_div/PartRem[44][3] ), .Y(
        \u_div/u_add_PartRem_2_43/n3 ) );
  OR2X2 U105 ( .A(\u_div/PartRem[37][2] ), .B(\u_div/PartRem[37][3] ), .Y(
        \u_div/u_add_PartRem_2_36/n3 ) );
  OR2X2 U106 ( .A(\u_div/PartRem[49][2] ), .B(\u_div/PartRem[49][3] ), .Y(
        \u_div/u_add_PartRem_2_48/n3 ) );
  OR2X2 U107 ( .A(\u_div/PartRem[46][2] ), .B(\u_div/PartRem[46][3] ), .Y(
        \u_div/u_add_PartRem_2_45/n3 ) );
  OR2X2 U108 ( .A(\u_div/PartRem[31][2] ), .B(\u_div/PartRem[31][3] ), .Y(
        \u_div/u_add_PartRem_2_30/n3 ) );
  OR2X2 U109 ( .A(\u_div/PartRem[40][2] ), .B(\u_div/PartRem[40][3] ), .Y(
        \u_div/u_add_PartRem_2_39/n3 ) );
  OR2X2 U110 ( .A(\u_div/PartRem[54][2] ), .B(\u_div/PartRem[54][3] ), .Y(
        \u_div/u_add_PartRem_2_53/n3 ) );
  OR2X2 U111 ( .A(\u_div/PartRem[47][2] ), .B(\u_div/PartRem[47][3] ), .Y(
        \u_div/u_add_PartRem_2_46/n3 ) );
  OR2X2 U112 ( .A(\u_div/PartRem[45][2] ), .B(\u_div/PartRem[45][3] ), .Y(
        \u_div/u_add_PartRem_2_44/n3 ) );
  OR2X2 U113 ( .A(\u_div/PartRem[50][2] ), .B(\u_div/PartRem[50][3] ), .Y(
        \u_div/u_add_PartRem_2_49/n3 ) );
  OR2X2 U114 ( .A(\u_div/PartRem[51][2] ), .B(\u_div/PartRem[51][3] ), .Y(
        \u_div/u_add_PartRem_2_50/n3 ) );
  OR2X2 U115 ( .A(\u_div/PartRem[57][2] ), .B(\u_div/PartRem[57][3] ), .Y(
        \u_div/u_add_PartRem_2_56/n3 ) );
  OR2X2 U116 ( .A(\u_div/PartRem[52][2] ), .B(\u_div/PartRem[52][3] ), .Y(
        \u_div/u_add_PartRem_2_51/n3 ) );
  OR2X2 U117 ( .A(\u_div/PartRem[55][2] ), .B(\u_div/PartRem[55][3] ), .Y(
        \u_div/u_add_PartRem_2_54/n3 ) );
  OR2X2 U118 ( .A(\u_div/PartRem[56][2] ), .B(\u_div/PartRem[56][3] ), .Y(
        \u_div/u_add_PartRem_2_55/n3 ) );
  OR2X2 U119 ( .A(\u_div/PartRem[58][2] ), .B(\u_div/PartRem[58][3] ), .Y(
        \u_div/u_add_PartRem_2_57/n3 ) );
  ADDHX2 U120 ( .A(\u_div/PartRem[59][4] ), .B(\u_div/u_add_PartRem_2_58/n3 ), 
        .CO(\u_div/u_add_PartRem_2_58/n2 ), .S(\u_div/SumTmp[58][4] ) );
  OR2X2 U121 ( .A(\u_div/PartRem[59][2] ), .B(\u_div/PartRem[59][3] ), .Y(
        \u_div/u_add_PartRem_2_58/n3 ) );
  OR2X2 U122 ( .A(\u_div/PartRem[15][2] ), .B(\u_div/PartRem[15][3] ), .Y(
        \u_div/u_add_PartRem_2_14/n3 ) );
  ADDHX1 U123 ( .A(\u_div/PartRem[4][4] ), .B(\u_div/u_add_PartRem_2_3/n3 ), 
        .CO(\u_div/u_add_PartRem_2_3/n2 ), .S(\u_div/SumTmp[3][4] ) );
  ADDHX1 U124 ( .A(\u_div/PartRem[2][4] ), .B(\u_div/u_add_PartRem_2_1/n3 ), 
        .CO(\u_div/u_add_PartRem_2_1/n2 ), .S(\u_div/SumTmp[1][4] ) );
  OR2X4 U125 ( .A(\u_div/PartRem[1][3] ), .B(\u_div/PartRem[1][2] ), .Y(n10)
         );
  ADDHX1 U126 ( .A(\u_div/PartRem[24][4] ), .B(\u_div/u_add_PartRem_2_23/n3 ), 
        .CO(\u_div/u_add_PartRem_2_23/n2 ), .S(\u_div/SumTmp[23][4] ) );
  ADDHX1 U127 ( .A(\u_div/PartRem[21][4] ), .B(\u_div/u_add_PartRem_2_20/n3 ), 
        .CO(\u_div/u_add_PartRem_2_20/n2 ), .S(\u_div/SumTmp[20][4] ) );
  ADDHX1 U128 ( .A(\u_div/PartRem[16][4] ), .B(\u_div/u_add_PartRem_2_15/n3 ), 
        .CO(\u_div/u_add_PartRem_2_15/n2 ), .S(\u_div/SumTmp[15][4] ) );
  ADDHX1 U129 ( .A(\u_div/PartRem[11][4] ), .B(\u_div/u_add_PartRem_2_10/n3 ), 
        .CO(\u_div/u_add_PartRem_2_10/n2 ), .S(\u_div/SumTmp[10][4] ) );
  ADDHX1 U130 ( .A(\u_div/PartRem[6][4] ), .B(\u_div/u_add_PartRem_2_5/n3 ), 
        .CO(\u_div/u_add_PartRem_2_5/n2 ), .S(\u_div/SumTmp[5][4] ) );
  OR2X1 U131 ( .A(\u_div/PartRem[53][2] ), .B(\u_div/PartRem[53][3] ), .Y(
        \u_div/u_add_PartRem_2_52/n3 ) );
  OR2X1 U132 ( .A(\u_div/PartRem[48][2] ), .B(\u_div/PartRem[48][3] ), .Y(
        \u_div/u_add_PartRem_2_47/n3 ) );
  OR2X1 U133 ( .A(\u_div/PartRem[43][2] ), .B(\u_div/PartRem[43][3] ), .Y(
        \u_div/u_add_PartRem_2_42/n3 ) );
  OR2X1 U134 ( .A(\u_div/PartRem[38][2] ), .B(\u_div/PartRem[38][3] ), .Y(
        \u_div/u_add_PartRem_2_37/n3 ) );
  OR2X1 U135 ( .A(\u_div/PartRem[33][2] ), .B(\u_div/PartRem[33][3] ), .Y(
        \u_div/u_add_PartRem_2_32/n3 ) );
  OR2X1 U136 ( .A(\u_div/PartRem[23][2] ), .B(\u_div/PartRem[23][3] ), .Y(
        \u_div/u_add_PartRem_2_22/n3 ) );
  OR2X1 U137 ( .A(\u_div/PartRem[18][2] ), .B(\u_div/PartRem[18][3] ), .Y(
        \u_div/u_add_PartRem_2_17/n3 ) );
  OR2X1 U138 ( .A(\u_div/PartRem[13][2] ), .B(\u_div/PartRem[13][3] ), .Y(
        \u_div/u_add_PartRem_2_12/n3 ) );
  OR2X1 U139 ( .A(\u_div/PartRem[8][2] ), .B(\u_div/PartRem[8][3] ), .Y(
        \u_div/u_add_PartRem_2_7/n3 ) );
  XNOR2XL U140 ( .A(\u_div/PartRem[64][0] ), .B(n12), .Y(\u_div/SumTmp[59][4] ) );
  XOR2XL U141 ( .A(\u_div/CryTmp[54][6] ), .B(n8), .Y(\u_div/QInv[54] ) );
  XOR2XL U142 ( .A(\u_div/CryTmp[52][6] ), .B(n9), .Y(\u_div/QInv[52] ) );
  XOR2XL U143 ( .A(\u_div/CryTmp[46][6] ), .B(n8), .Y(\u_div/QInv[46] ) );
  XOR2XL U144 ( .A(\u_div/CryTmp[44][6] ), .B(n9), .Y(\u_div/QInv[44] ) );
  XOR2XL U145 ( .A(\u_div/CryTmp[35][6] ), .B(n8), .Y(\u_div/QInv[35] ) );
  XOR2XL U146 ( .A(\u_div/CryTmp[34][6] ), .B(n9), .Y(\u_div/QInv[34] ) );
  XOR2XL U147 ( .A(\u_div/CryTmp[36][6] ), .B(n9), .Y(\u_div/QInv[36] ) );
  XOR2XL U148 ( .A(\u_div/CryTmp[26][6] ), .B(n9), .Y(\u_div/QInv[26] ) );
  XOR2XL U149 ( .A(\u_div/CryTmp[25][6] ), .B(n8), .Y(\u_div/QInv[25] ) );
  XOR2XL U150 ( .A(\u_div/CryTmp[16][6] ), .B(n9), .Y(\u_div/QInv[16] ) );
  XOR2XL U151 ( .A(\u_div/CryTmp[15][6] ), .B(n8), .Y(\u_div/QInv[15] ) );
  XOR2XL U152 ( .A(\u_div/CryTmp[14][6] ), .B(n9), .Y(\u_div/QInv[14] ) );
  XOR2XL U153 ( .A(\u_div/CryTmp[5][6] ), .B(n8), .Y(\u_div/QInv[5] ) );
  XOR2XL U154 ( .A(\u_div/CryTmp[6][6] ), .B(n9), .Y(\u_div/QInv[6] ) );
  XOR2XL U155 ( .A(\u_div/CryTmp[53][6] ), .B(n7), .Y(\u_div/QInv[53] ) );
  XOR2XL U156 ( .A(\u_div/CryTmp[45][6] ), .B(n7), .Y(\u_div/QInv[45] ) );
  XOR2XL U157 ( .A(\u_div/CryTmp[24][6] ), .B(n7), .Y(\u_div/QInv[24] ) );
  INVXL U158 ( .A(\u_div/PartRem[23][2] ), .Y(\u_div/SumTmp[22][2] ) );
  INVXL U159 ( .A(\u_div/PartRem[18][2] ), .Y(\u_div/SumTmp[17][2] ) );
  INVXL U160 ( .A(\u_div/PartRem[13][2] ), .Y(\u_div/SumTmp[12][2] ) );
  INVXL U161 ( .A(\u_div/PartRem[8][2] ), .Y(\u_div/SumTmp[7][2] ) );
  INVXL U162 ( .A(\u_div/PartRem[59][2] ), .Y(\u_div/SumTmp[58][2] ) );
  INVX3 U163 ( .A(n6), .Y(n7) );
  INVXL U164 ( .A(\u_div/PartRem[2][2] ), .Y(\u_div/SumTmp[1][2] ) );
  CLKINVX1 U165 ( .A(\u_div/QInv[63] ), .Y(n6) );
  OR2X2 U166 ( .A(\u_div/PartRem[3][5] ), .B(\u_div/u_add_PartRem_2_2/n2 ), 
        .Y(\u_div/CryTmp[2][6] ) );
  OR2X1 U167 ( .A(\u_div/PartRem[2][5] ), .B(\u_div/u_add_PartRem_2_1/n2 ), 
        .Y(\u_div/CryTmp[1][6] ) );
  XOR2X1 U168 ( .A(\u_div/CryTmp[0][6] ), .B(n9), .Y(\u_div/QInv[0] ) );
  AO21X1 U169 ( .A0(\u_div/PartRem[1][4] ), .A1(n10), .B0(
        \u_div/PartRem[1][5] ), .Y(\u_div/CryTmp[0][6] ) );
  OR2X1 U170 ( .A(\u_div/PartRem[28][2] ), .B(\u_div/PartRem[28][3] ), .Y(
        \u_div/u_add_PartRem_2_27/n3 ) );
  MXI2X1 U171 ( .A(n11), .B(\u_div/PartRem[62][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(\u_div/PartRem[59][3] ) );
  CLKINVX1 U172 ( .A(\u_div/PartRem[62][0] ), .Y(n11) );
  MXI2X1 U173 ( .A(\u_div/SumTmp[58][2] ), .B(\u_div/PartRem[59][2] ), .S0(
        \u_div/CryTmp[58][6] ), .Y(\u_div/PartRem[58][3] ) );
  MXI2X1 U174 ( .A(\u_div/SumTmp[57][2] ), .B(\u_div/PartRem[58][2] ), .S0(
        \u_div/CryTmp[57][6] ), .Y(\u_div/PartRem[57][3] ) );
  CLKINVX1 U175 ( .A(\u_div/PartRem[58][2] ), .Y(\u_div/SumTmp[57][2] ) );
  MXI2X1 U176 ( .A(\u_div/SumTmp[56][2] ), .B(\u_div/PartRem[57][2] ), .S0(
        \u_div/CryTmp[56][6] ), .Y(\u_div/PartRem[56][3] ) );
  CLKINVX1 U177 ( .A(\u_div/PartRem[57][2] ), .Y(\u_div/SumTmp[56][2] ) );
  MXI2X1 U178 ( .A(\u_div/SumTmp[54][2] ), .B(\u_div/PartRem[55][2] ), .S0(
        \u_div/CryTmp[54][6] ), .Y(\u_div/PartRem[54][3] ) );
  CLKINVX1 U179 ( .A(\u_div/PartRem[55][2] ), .Y(\u_div/SumTmp[54][2] ) );
  MXI2X1 U180 ( .A(\u_div/SumTmp[55][2] ), .B(\u_div/PartRem[56][2] ), .S0(
        \u_div/CryTmp[55][6] ), .Y(\u_div/PartRem[55][3] ) );
  CLKINVX1 U181 ( .A(\u_div/PartRem[56][2] ), .Y(\u_div/SumTmp[55][2] ) );
  MXI2X1 U182 ( .A(\u_div/SumTmp[52][2] ), .B(\u_div/PartRem[53][2] ), .S0(
        \u_div/CryTmp[52][6] ), .Y(\u_div/PartRem[52][3] ) );
  CLKINVX1 U183 ( .A(\u_div/PartRem[53][2] ), .Y(\u_div/SumTmp[52][2] ) );
  MXI2X1 U184 ( .A(\u_div/SumTmp[51][2] ), .B(\u_div/PartRem[52][2] ), .S0(
        \u_div/CryTmp[51][6] ), .Y(\u_div/PartRem[51][3] ) );
  CLKINVX1 U185 ( .A(\u_div/PartRem[52][2] ), .Y(\u_div/SumTmp[51][2] ) );
  MXI2X1 U186 ( .A(\u_div/SumTmp[49][2] ), .B(\u_div/PartRem[50][2] ), .S0(
        \u_div/CryTmp[49][6] ), .Y(\u_div/PartRem[49][3] ) );
  CLKINVX1 U187 ( .A(\u_div/PartRem[50][2] ), .Y(\u_div/SumTmp[49][2] ) );
  MXI2X1 U188 ( .A(\u_div/SumTmp[50][2] ), .B(\u_div/PartRem[51][2] ), .S0(
        \u_div/CryTmp[50][6] ), .Y(\u_div/PartRem[50][3] ) );
  CLKINVX1 U189 ( .A(\u_div/PartRem[51][2] ), .Y(\u_div/SumTmp[50][2] ) );
  MXI2X1 U190 ( .A(\u_div/SumTmp[47][2] ), .B(\u_div/PartRem[48][2] ), .S0(
        \u_div/CryTmp[47][6] ), .Y(\u_div/PartRem[47][3] ) );
  CLKINVX1 U191 ( .A(\u_div/PartRem[48][2] ), .Y(\u_div/SumTmp[47][2] ) );
  MXI2X1 U192 ( .A(\u_div/SumTmp[46][2] ), .B(\u_div/PartRem[47][2] ), .S0(
        \u_div/CryTmp[46][6] ), .Y(\u_div/PartRem[46][3] ) );
  CLKINVX1 U193 ( .A(\u_div/PartRem[47][2] ), .Y(\u_div/SumTmp[46][2] ) );
  MXI2X1 U194 ( .A(\u_div/SumTmp[44][2] ), .B(\u_div/PartRem[45][2] ), .S0(
        \u_div/CryTmp[44][6] ), .Y(\u_div/PartRem[44][3] ) );
  CLKINVX1 U195 ( .A(\u_div/PartRem[45][2] ), .Y(\u_div/SumTmp[44][2] ) );
  MXI2X1 U196 ( .A(\u_div/SumTmp[45][2] ), .B(\u_div/PartRem[46][2] ), .S0(
        \u_div/CryTmp[45][6] ), .Y(\u_div/PartRem[45][3] ) );
  CLKINVX1 U197 ( .A(\u_div/PartRem[46][2] ), .Y(\u_div/SumTmp[45][2] ) );
  MXI2X1 U198 ( .A(\u_div/SumTmp[42][2] ), .B(\u_div/PartRem[43][2] ), .S0(
        \u_div/CryTmp[42][6] ), .Y(\u_div/PartRem[42][3] ) );
  CLKINVX1 U199 ( .A(\u_div/PartRem[43][2] ), .Y(\u_div/SumTmp[42][2] ) );
  MXI2X1 U200 ( .A(\u_div/SumTmp[41][2] ), .B(\u_div/PartRem[42][2] ), .S0(
        \u_div/CryTmp[41][6] ), .Y(\u_div/PartRem[41][3] ) );
  CLKINVX1 U201 ( .A(\u_div/PartRem[42][2] ), .Y(\u_div/SumTmp[41][2] ) );
  MXI2X1 U202 ( .A(\u_div/SumTmp[39][2] ), .B(\u_div/PartRem[40][2] ), .S0(
        \u_div/CryTmp[39][6] ), .Y(\u_div/PartRem[39][3] ) );
  CLKINVX1 U203 ( .A(\u_div/PartRem[40][2] ), .Y(\u_div/SumTmp[39][2] ) );
  MXI2X1 U204 ( .A(\u_div/SumTmp[40][2] ), .B(\u_div/PartRem[41][2] ), .S0(
        \u_div/CryTmp[40][6] ), .Y(\u_div/PartRem[40][3] ) );
  CLKINVX1 U205 ( .A(\u_div/PartRem[41][2] ), .Y(\u_div/SumTmp[40][2] ) );
  MXI2X1 U206 ( .A(\u_div/SumTmp[37][2] ), .B(\u_div/PartRem[38][2] ), .S0(
        \u_div/CryTmp[37][6] ), .Y(\u_div/PartRem[37][3] ) );
  CLKINVX1 U207 ( .A(\u_div/PartRem[38][2] ), .Y(\u_div/SumTmp[37][2] ) );
  MXI2X1 U208 ( .A(\u_div/SumTmp[36][2] ), .B(\u_div/PartRem[37][2] ), .S0(
        \u_div/CryTmp[36][6] ), .Y(\u_div/PartRem[36][3] ) );
  CLKINVX1 U209 ( .A(\u_div/PartRem[37][2] ), .Y(\u_div/SumTmp[36][2] ) );
  MXI2X1 U210 ( .A(\u_div/SumTmp[34][2] ), .B(\u_div/PartRem[35][2] ), .S0(
        \u_div/CryTmp[34][6] ), .Y(\u_div/PartRem[34][3] ) );
  CLKINVX1 U211 ( .A(\u_div/PartRem[35][2] ), .Y(\u_div/SumTmp[34][2] ) );
  MXI2X1 U212 ( .A(\u_div/SumTmp[35][2] ), .B(\u_div/PartRem[36][2] ), .S0(
        \u_div/CryTmp[35][6] ), .Y(\u_div/PartRem[35][3] ) );
  CLKINVX1 U213 ( .A(\u_div/PartRem[36][2] ), .Y(\u_div/SumTmp[35][2] ) );
  MXI2X1 U214 ( .A(\u_div/SumTmp[32][2] ), .B(\u_div/PartRem[33][2] ), .S0(
        \u_div/CryTmp[32][6] ), .Y(\u_div/PartRem[32][3] ) );
  CLKINVX1 U215 ( .A(\u_div/PartRem[33][2] ), .Y(\u_div/SumTmp[32][2] ) );
  MXI2X1 U216 ( .A(\u_div/SumTmp[31][2] ), .B(\u_div/PartRem[32][2] ), .S0(
        \u_div/CryTmp[31][6] ), .Y(\u_div/PartRem[31][3] ) );
  CLKINVX1 U217 ( .A(\u_div/PartRem[32][2] ), .Y(\u_div/SumTmp[31][2] ) );
  MXI2X1 U218 ( .A(\u_div/SumTmp[29][2] ), .B(\u_div/PartRem[30][2] ), .S0(
        \u_div/CryTmp[29][6] ), .Y(\u_div/PartRem[29][3] ) );
  CLKINVX1 U219 ( .A(\u_div/PartRem[30][2] ), .Y(\u_div/SumTmp[29][2] ) );
  MXI2X1 U220 ( .A(\u_div/SumTmp[30][2] ), .B(\u_div/PartRem[31][2] ), .S0(
        \u_div/CryTmp[30][6] ), .Y(\u_div/PartRem[30][3] ) );
  CLKINVX1 U221 ( .A(\u_div/PartRem[31][2] ), .Y(\u_div/SumTmp[30][2] ) );
  MXI2X1 U222 ( .A(\u_div/SumTmp[27][2] ), .B(\u_div/PartRem[28][2] ), .S0(
        \u_div/CryTmp[27][6] ), .Y(\u_div/PartRem[27][3] ) );
  CLKINVX1 U223 ( .A(\u_div/PartRem[28][2] ), .Y(\u_div/SumTmp[27][2] ) );
  MXI2X1 U224 ( .A(\u_div/SumTmp[26][2] ), .B(\u_div/PartRem[27][2] ), .S0(
        \u_div/CryTmp[26][6] ), .Y(\u_div/PartRem[26][3] ) );
  CLKINVX1 U225 ( .A(\u_div/PartRem[27][2] ), .Y(\u_div/SumTmp[26][2] ) );
  MXI2X1 U226 ( .A(\u_div/SumTmp[25][2] ), .B(\u_div/PartRem[26][2] ), .S0(
        \u_div/CryTmp[25][6] ), .Y(\u_div/PartRem[25][3] ) );
  CLKINVX1 U227 ( .A(\u_div/PartRem[26][2] ), .Y(\u_div/SumTmp[25][2] ) );
  CLKINVX1 U228 ( .A(\u_div/PartRem[25][2] ), .Y(\u_div/SumTmp[24][2] ) );
  MXI2X1 U229 ( .A(\u_div/SumTmp[22][2] ), .B(\u_div/PartRem[23][2] ), .S0(
        \u_div/CryTmp[22][6] ), .Y(\u_div/PartRem[22][3] ) );
  CLKINVX1 U230 ( .A(\u_div/PartRem[22][2] ), .Y(\u_div/SumTmp[21][2] ) );
  MXI2X1 U231 ( .A(\u_div/SumTmp[17][2] ), .B(\u_div/PartRem[18][2] ), .S0(
        \u_div/CryTmp[17][6] ), .Y(\u_div/PartRem[17][3] ) );
  CLKINVX1 U232 ( .A(\u_div/PartRem[17][2] ), .Y(\u_div/SumTmp[16][2] ) );
  MXI2X1 U233 ( .A(\u_div/SumTmp[12][2] ), .B(\u_div/PartRem[13][2] ), .S0(
        \u_div/CryTmp[12][6] ), .Y(\u_div/PartRem[12][3] ) );
  CLKINVX1 U234 ( .A(\u_div/PartRem[12][2] ), .Y(\u_div/SumTmp[11][2] ) );
  MXI2X1 U235 ( .A(\u_div/SumTmp[7][2] ), .B(\u_div/PartRem[8][2] ), .S0(
        \u_div/CryTmp[7][6] ), .Y(\u_div/PartRem[7][3] ) );
  CLKINVX1 U236 ( .A(\u_div/PartRem[7][2] ), .Y(\u_div/SumTmp[6][2] ) );
  MXI2X1 U237 ( .A(\u_div/SumTmp[3][2] ), .B(\u_div/PartRem[4][2] ), .S0(
        \u_div/CryTmp[3][6] ), .Y(\u_div/PartRem[3][3] ) );
  CLKINVX1 U238 ( .A(\u_div/PartRem[4][2] ), .Y(\u_div/SumTmp[3][2] ) );
  MXI2X1 U239 ( .A(\u_div/SumTmp[23][2] ), .B(\u_div/PartRem[24][2] ), .S0(
        \u_div/CryTmp[23][6] ), .Y(\u_div/PartRem[23][3] ) );
  CLKINVX1 U240 ( .A(\u_div/PartRem[24][2] ), .Y(\u_div/SumTmp[23][2] ) );
  MXI2X1 U241 ( .A(\u_div/SumTmp[18][2] ), .B(\u_div/PartRem[19][2] ), .S0(
        \u_div/CryTmp[18][6] ), .Y(\u_div/PartRem[18][3] ) );
  CLKINVX1 U242 ( .A(\u_div/PartRem[19][2] ), .Y(\u_div/SumTmp[18][2] ) );
  MXI2X1 U243 ( .A(\u_div/SumTmp[13][2] ), .B(\u_div/PartRem[14][2] ), .S0(
        \u_div/CryTmp[13][6] ), .Y(\u_div/PartRem[13][3] ) );
  CLKINVX1 U244 ( .A(\u_div/PartRem[14][2] ), .Y(\u_div/SumTmp[13][2] ) );
  MXI2X1 U245 ( .A(\u_div/SumTmp[8][2] ), .B(\u_div/PartRem[9][2] ), .S0(
        \u_div/CryTmp[8][6] ), .Y(\u_div/PartRem[8][3] ) );
  CLKINVX1 U246 ( .A(\u_div/PartRem[9][2] ), .Y(\u_div/SumTmp[8][2] ) );
  MXI2X1 U247 ( .A(\u_div/SumTmp[20][2] ), .B(\u_div/PartRem[21][2] ), .S0(
        \u_div/CryTmp[20][6] ), .Y(\u_div/PartRem[20][3] ) );
  CLKINVX1 U248 ( .A(\u_div/PartRem[21][2] ), .Y(\u_div/SumTmp[20][2] ) );
  MXI2X1 U249 ( .A(\u_div/SumTmp[15][2] ), .B(\u_div/PartRem[16][2] ), .S0(
        \u_div/CryTmp[15][6] ), .Y(\u_div/PartRem[15][3] ) );
  CLKINVX1 U250 ( .A(\u_div/PartRem[16][2] ), .Y(\u_div/SumTmp[15][2] ) );
  MXI2X1 U251 ( .A(\u_div/SumTmp[10][2] ), .B(\u_div/PartRem[11][2] ), .S0(
        \u_div/CryTmp[10][6] ), .Y(\u_div/PartRem[10][3] ) );
  CLKINVX1 U252 ( .A(\u_div/PartRem[11][2] ), .Y(\u_div/SumTmp[10][2] ) );
  MXI2X1 U253 ( .A(\u_div/SumTmp[5][2] ), .B(\u_div/PartRem[6][2] ), .S0(
        \u_div/CryTmp[5][6] ), .Y(\u_div/PartRem[5][3] ) );
  CLKINVX1 U254 ( .A(\u_div/PartRem[6][2] ), .Y(\u_div/SumTmp[5][2] ) );
  MXI2X1 U255 ( .A(\u_div/SumTmp[53][2] ), .B(\u_div/PartRem[54][2] ), .S0(
        \u_div/CryTmp[53][6] ), .Y(\u_div/PartRem[53][3] ) );
  CLKINVX1 U256 ( .A(\u_div/PartRem[54][2] ), .Y(\u_div/SumTmp[53][2] ) );
  MXI2X1 U257 ( .A(\u_div/SumTmp[48][2] ), .B(\u_div/PartRem[49][2] ), .S0(
        \u_div/CryTmp[48][6] ), .Y(\u_div/PartRem[48][3] ) );
  CLKINVX1 U258 ( .A(\u_div/PartRem[49][2] ), .Y(\u_div/SumTmp[48][2] ) );
  MXI2X1 U259 ( .A(\u_div/SumTmp[43][2] ), .B(\u_div/PartRem[44][2] ), .S0(
        \u_div/CryTmp[43][6] ), .Y(\u_div/PartRem[43][3] ) );
  CLKINVX1 U260 ( .A(\u_div/PartRem[44][2] ), .Y(\u_div/SumTmp[43][2] ) );
  MXI2X1 U261 ( .A(\u_div/SumTmp[38][2] ), .B(\u_div/PartRem[39][2] ), .S0(
        \u_div/CryTmp[38][6] ), .Y(\u_div/PartRem[38][3] ) );
  CLKINVX1 U262 ( .A(\u_div/PartRem[39][2] ), .Y(\u_div/SumTmp[38][2] ) );
  MXI2X1 U263 ( .A(\u_div/SumTmp[33][2] ), .B(\u_div/PartRem[34][2] ), .S0(
        \u_div/CryTmp[33][6] ), .Y(\u_div/PartRem[33][3] ) );
  CLKINVX1 U264 ( .A(\u_div/PartRem[34][2] ), .Y(\u_div/SumTmp[33][2] ) );
  CLKINVX1 U265 ( .A(\u_div/PartRem[29][2] ), .Y(\u_div/SumTmp[28][2] ) );
  INVX4 U266 ( .A(n6), .Y(n9) );
  INVX4 U267 ( .A(n6), .Y(n8) );
  OR2X1 U268 ( .A(\u_div/PartRem[59][5] ), .B(\u_div/u_add_PartRem_2_58/n2 ), 
        .Y(\u_div/CryTmp[58][6] ) );
  XNOR2X1 U269 ( .A(\u_div/PartRem[59][3] ), .B(\u_div/PartRem[59][2] ), .Y(
        \u_div/SumTmp[58][3] ) );
  OR2X1 U270 ( .A(\u_div/PartRem[58][5] ), .B(\u_div/u_add_PartRem_2_57/n2 ), 
        .Y(\u_div/CryTmp[57][6] ) );
  XNOR2X1 U271 ( .A(\u_div/PartRem[58][3] ), .B(\u_div/PartRem[58][2] ), .Y(
        \u_div/SumTmp[57][3] ) );
  OR2X1 U272 ( .A(\u_div/PartRem[57][5] ), .B(\u_div/u_add_PartRem_2_56/n2 ), 
        .Y(\u_div/CryTmp[56][6] ) );
  XNOR2X1 U273 ( .A(\u_div/PartRem[57][3] ), .B(\u_div/PartRem[57][2] ), .Y(
        \u_div/SumTmp[56][3] ) );
  OR2X1 U274 ( .A(\u_div/PartRem[56][5] ), .B(\u_div/u_add_PartRem_2_55/n2 ), 
        .Y(\u_div/CryTmp[55][6] ) );
  XNOR2X1 U275 ( .A(\u_div/PartRem[56][3] ), .B(\u_div/PartRem[56][2] ), .Y(
        \u_div/SumTmp[55][3] ) );
  OR2X1 U276 ( .A(\u_div/PartRem[55][5] ), .B(\u_div/u_add_PartRem_2_54/n2 ), 
        .Y(\u_div/CryTmp[54][6] ) );
  XNOR2X1 U277 ( .A(\u_div/PartRem[55][3] ), .B(\u_div/PartRem[55][2] ), .Y(
        \u_div/SumTmp[54][3] ) );
  OR2X1 U278 ( .A(\u_div/PartRem[54][5] ), .B(\u_div/u_add_PartRem_2_53/n2 ), 
        .Y(\u_div/CryTmp[53][6] ) );
  XNOR2X1 U279 ( .A(\u_div/PartRem[54][3] ), .B(\u_div/PartRem[54][2] ), .Y(
        \u_div/SumTmp[53][3] ) );
  OR2X1 U280 ( .A(\u_div/PartRem[53][5] ), .B(\u_div/u_add_PartRem_2_52/n2 ), 
        .Y(\u_div/CryTmp[52][6] ) );
  XNOR2X1 U281 ( .A(\u_div/PartRem[53][3] ), .B(\u_div/PartRem[53][2] ), .Y(
        \u_div/SumTmp[52][3] ) );
  OR2X1 U282 ( .A(\u_div/PartRem[52][5] ), .B(\u_div/u_add_PartRem_2_51/n2 ), 
        .Y(\u_div/CryTmp[51][6] ) );
  XNOR2X1 U283 ( .A(\u_div/PartRem[52][3] ), .B(\u_div/PartRem[52][2] ), .Y(
        \u_div/SumTmp[51][3] ) );
  OR2X1 U284 ( .A(\u_div/PartRem[51][5] ), .B(\u_div/u_add_PartRem_2_50/n2 ), 
        .Y(\u_div/CryTmp[50][6] ) );
  XNOR2X1 U285 ( .A(\u_div/PartRem[51][3] ), .B(\u_div/PartRem[51][2] ), .Y(
        \u_div/SumTmp[50][3] ) );
  OR2X1 U286 ( .A(\u_div/PartRem[50][5] ), .B(\u_div/u_add_PartRem_2_49/n2 ), 
        .Y(\u_div/CryTmp[49][6] ) );
  XNOR2X1 U287 ( .A(\u_div/PartRem[50][3] ), .B(\u_div/PartRem[50][2] ), .Y(
        \u_div/SumTmp[49][3] ) );
  OR2X1 U288 ( .A(\u_div/PartRem[49][5] ), .B(\u_div/u_add_PartRem_2_48/n2 ), 
        .Y(\u_div/CryTmp[48][6] ) );
  XNOR2X1 U289 ( .A(\u_div/PartRem[49][3] ), .B(\u_div/PartRem[49][2] ), .Y(
        \u_div/SumTmp[48][3] ) );
  OR2X1 U290 ( .A(\u_div/PartRem[48][5] ), .B(\u_div/u_add_PartRem_2_47/n2 ), 
        .Y(\u_div/CryTmp[47][6] ) );
  XNOR2X1 U291 ( .A(\u_div/PartRem[48][3] ), .B(\u_div/PartRem[48][2] ), .Y(
        \u_div/SumTmp[47][3] ) );
  OR2X1 U292 ( .A(\u_div/PartRem[47][5] ), .B(\u_div/u_add_PartRem_2_46/n2 ), 
        .Y(\u_div/CryTmp[46][6] ) );
  XNOR2X1 U293 ( .A(\u_div/PartRem[47][3] ), .B(\u_div/PartRem[47][2] ), .Y(
        \u_div/SumTmp[46][3] ) );
  OR2X1 U294 ( .A(\u_div/PartRem[46][5] ), .B(\u_div/u_add_PartRem_2_45/n2 ), 
        .Y(\u_div/CryTmp[45][6] ) );
  XNOR2X1 U295 ( .A(\u_div/PartRem[46][3] ), .B(\u_div/PartRem[46][2] ), .Y(
        \u_div/SumTmp[45][3] ) );
  OR2X1 U296 ( .A(\u_div/PartRem[45][5] ), .B(\u_div/u_add_PartRem_2_44/n2 ), 
        .Y(\u_div/CryTmp[44][6] ) );
  XNOR2X1 U297 ( .A(\u_div/PartRem[45][3] ), .B(\u_div/PartRem[45][2] ), .Y(
        \u_div/SumTmp[44][3] ) );
  OR2X1 U298 ( .A(\u_div/PartRem[44][5] ), .B(\u_div/u_add_PartRem_2_43/n2 ), 
        .Y(\u_div/CryTmp[43][6] ) );
  XNOR2X1 U299 ( .A(\u_div/PartRem[44][3] ), .B(\u_div/PartRem[44][2] ), .Y(
        \u_div/SumTmp[43][3] ) );
  OR2X1 U300 ( .A(\u_div/PartRem[43][5] ), .B(\u_div/u_add_PartRem_2_42/n2 ), 
        .Y(\u_div/CryTmp[42][6] ) );
  XNOR2X1 U301 ( .A(\u_div/PartRem[43][3] ), .B(\u_div/PartRem[43][2] ), .Y(
        \u_div/SumTmp[42][3] ) );
  OR2X1 U302 ( .A(\u_div/PartRem[42][5] ), .B(\u_div/u_add_PartRem_2_41/n2 ), 
        .Y(\u_div/CryTmp[41][6] ) );
  XNOR2X1 U303 ( .A(\u_div/PartRem[42][3] ), .B(\u_div/PartRem[42][2] ), .Y(
        \u_div/SumTmp[41][3] ) );
  OR2X1 U304 ( .A(\u_div/PartRem[41][5] ), .B(\u_div/u_add_PartRem_2_40/n2 ), 
        .Y(\u_div/CryTmp[40][6] ) );
  XNOR2X1 U305 ( .A(\u_div/PartRem[41][3] ), .B(\u_div/PartRem[41][2] ), .Y(
        \u_div/SumTmp[40][3] ) );
  OR2X1 U306 ( .A(\u_div/PartRem[40][5] ), .B(\u_div/u_add_PartRem_2_39/n2 ), 
        .Y(\u_div/CryTmp[39][6] ) );
  XNOR2X1 U307 ( .A(\u_div/PartRem[40][3] ), .B(\u_div/PartRem[40][2] ), .Y(
        \u_div/SumTmp[39][3] ) );
  OR2X1 U308 ( .A(\u_div/PartRem[39][5] ), .B(\u_div/u_add_PartRem_2_38/n2 ), 
        .Y(\u_div/CryTmp[38][6] ) );
  XNOR2X1 U309 ( .A(\u_div/PartRem[39][3] ), .B(\u_div/PartRem[39][2] ), .Y(
        \u_div/SumTmp[38][3] ) );
  OR2X1 U310 ( .A(\u_div/PartRem[38][5] ), .B(\u_div/u_add_PartRem_2_37/n2 ), 
        .Y(\u_div/CryTmp[37][6] ) );
  XNOR2X1 U311 ( .A(\u_div/PartRem[38][3] ), .B(\u_div/PartRem[38][2] ), .Y(
        \u_div/SumTmp[37][3] ) );
  OR2X1 U312 ( .A(\u_div/PartRem[37][5] ), .B(\u_div/u_add_PartRem_2_36/n2 ), 
        .Y(\u_div/CryTmp[36][6] ) );
  XNOR2X1 U313 ( .A(\u_div/PartRem[37][3] ), .B(\u_div/PartRem[37][2] ), .Y(
        \u_div/SumTmp[36][3] ) );
  OR2X1 U314 ( .A(\u_div/PartRem[36][5] ), .B(\u_div/u_add_PartRem_2_35/n2 ), 
        .Y(\u_div/CryTmp[35][6] ) );
  XNOR2X1 U315 ( .A(\u_div/PartRem[36][3] ), .B(\u_div/PartRem[36][2] ), .Y(
        \u_div/SumTmp[35][3] ) );
  OR2X1 U316 ( .A(\u_div/PartRem[35][5] ), .B(\u_div/u_add_PartRem_2_34/n2 ), 
        .Y(\u_div/CryTmp[34][6] ) );
  XNOR2X1 U317 ( .A(\u_div/PartRem[35][3] ), .B(\u_div/PartRem[35][2] ), .Y(
        \u_div/SumTmp[34][3] ) );
  OR2X1 U318 ( .A(\u_div/PartRem[34][5] ), .B(\u_div/u_add_PartRem_2_33/n2 ), 
        .Y(\u_div/CryTmp[33][6] ) );
  XNOR2X1 U319 ( .A(\u_div/PartRem[34][3] ), .B(\u_div/PartRem[34][2] ), .Y(
        \u_div/SumTmp[33][3] ) );
  OR2X1 U320 ( .A(\u_div/PartRem[33][5] ), .B(\u_div/u_add_PartRem_2_32/n2 ), 
        .Y(\u_div/CryTmp[32][6] ) );
  XNOR2X1 U321 ( .A(\u_div/PartRem[33][3] ), .B(\u_div/PartRem[33][2] ), .Y(
        \u_div/SumTmp[32][3] ) );
  OR2X1 U322 ( .A(\u_div/PartRem[32][5] ), .B(\u_div/u_add_PartRem_2_31/n2 ), 
        .Y(\u_div/CryTmp[31][6] ) );
  XNOR2X1 U323 ( .A(\u_div/PartRem[32][3] ), .B(\u_div/PartRem[32][2] ), .Y(
        \u_div/SumTmp[31][3] ) );
  OR2X1 U324 ( .A(\u_div/PartRem[31][5] ), .B(\u_div/u_add_PartRem_2_30/n2 ), 
        .Y(\u_div/CryTmp[30][6] ) );
  XNOR2X1 U325 ( .A(\u_div/PartRem[31][3] ), .B(\u_div/PartRem[31][2] ), .Y(
        \u_div/SumTmp[30][3] ) );
  OR2X1 U326 ( .A(\u_div/PartRem[30][5] ), .B(\u_div/u_add_PartRem_2_29/n2 ), 
        .Y(\u_div/CryTmp[29][6] ) );
  XNOR2X1 U327 ( .A(\u_div/PartRem[30][3] ), .B(\u_div/PartRem[30][2] ), .Y(
        \u_div/SumTmp[29][3] ) );
  OR2X1 U328 ( .A(\u_div/PartRem[29][5] ), .B(\u_div/u_add_PartRem_2_28/n2 ), 
        .Y(\u_div/CryTmp[28][6] ) );
  XNOR2X1 U329 ( .A(\u_div/PartRem[29][3] ), .B(\u_div/PartRem[29][2] ), .Y(
        \u_div/SumTmp[28][3] ) );
  OR2X1 U330 ( .A(\u_div/PartRem[28][5] ), .B(\u_div/u_add_PartRem_2_27/n2 ), 
        .Y(\u_div/CryTmp[27][6] ) );
  XNOR2X1 U331 ( .A(\u_div/PartRem[28][3] ), .B(\u_div/PartRem[28][2] ), .Y(
        \u_div/SumTmp[27][3] ) );
  OR2X1 U332 ( .A(\u_div/PartRem[27][5] ), .B(\u_div/u_add_PartRem_2_26/n2 ), 
        .Y(\u_div/CryTmp[26][6] ) );
  XNOR2X1 U333 ( .A(\u_div/PartRem[27][3] ), .B(\u_div/PartRem[27][2] ), .Y(
        \u_div/SumTmp[26][3] ) );
  OR2X1 U334 ( .A(\u_div/PartRem[26][5] ), .B(\u_div/u_add_PartRem_2_25/n2 ), 
        .Y(\u_div/CryTmp[25][6] ) );
  XNOR2X1 U335 ( .A(\u_div/PartRem[26][3] ), .B(\u_div/PartRem[26][2] ), .Y(
        \u_div/SumTmp[25][3] ) );
  OR2X1 U336 ( .A(\u_div/PartRem[25][5] ), .B(\u_div/u_add_PartRem_2_24/n2 ), 
        .Y(\u_div/CryTmp[24][6] ) );
  XNOR2X1 U337 ( .A(\u_div/PartRem[25][3] ), .B(\u_div/PartRem[25][2] ), .Y(
        \u_div/SumTmp[24][3] ) );
  XNOR2X1 U338 ( .A(\u_div/PartRem[24][3] ), .B(\u_div/PartRem[24][2] ), .Y(
        \u_div/SumTmp[23][3] ) );
  OR2X1 U339 ( .A(\u_div/PartRem[24][2] ), .B(\u_div/PartRem[24][3] ), .Y(
        \u_div/u_add_PartRem_2_23/n3 ) );
  OR2X1 U340 ( .A(\u_div/PartRem[23][5] ), .B(\u_div/u_add_PartRem_2_22/n2 ), 
        .Y(\u_div/CryTmp[22][6] ) );
  XNOR2X1 U341 ( .A(\u_div/PartRem[23][3] ), .B(\u_div/PartRem[23][2] ), .Y(
        \u_div/SumTmp[22][3] ) );
  XNOR2X1 U342 ( .A(\u_div/PartRem[22][3] ), .B(\u_div/PartRem[22][2] ), .Y(
        \u_div/SumTmp[21][3] ) );
  XNOR2X1 U343 ( .A(\u_div/PartRem[21][3] ), .B(\u_div/PartRem[21][2] ), .Y(
        \u_div/SumTmp[20][3] ) );
  OR2X1 U344 ( .A(\u_div/PartRem[21][2] ), .B(\u_div/PartRem[21][3] ), .Y(
        \u_div/u_add_PartRem_2_20/n3 ) );
  XNOR2X1 U345 ( .A(\u_div/PartRem[20][3] ), .B(\u_div/PartRem[20][2] ), .Y(
        \u_div/SumTmp[19][3] ) );
  XNOR2X1 U346 ( .A(\u_div/PartRem[19][3] ), .B(\u_div/PartRem[19][2] ), .Y(
        \u_div/SumTmp[18][3] ) );
  OR2X1 U347 ( .A(\u_div/PartRem[19][2] ), .B(\u_div/PartRem[19][3] ), .Y(
        \u_div/u_add_PartRem_2_18/n3 ) );
  OR2X1 U348 ( .A(\u_div/PartRem[18][5] ), .B(\u_div/u_add_PartRem_2_17/n2 ), 
        .Y(\u_div/CryTmp[17][6] ) );
  XNOR2X1 U349 ( .A(\u_div/PartRem[18][3] ), .B(\u_div/PartRem[18][2] ), .Y(
        \u_div/SumTmp[17][3] ) );
  XNOR2X1 U350 ( .A(\u_div/PartRem[17][3] ), .B(\u_div/PartRem[17][2] ), .Y(
        \u_div/SumTmp[16][3] ) );
  XNOR2X1 U351 ( .A(\u_div/PartRem[16][3] ), .B(\u_div/PartRem[16][2] ), .Y(
        \u_div/SumTmp[15][3] ) );
  OR2X1 U352 ( .A(\u_div/PartRem[16][2] ), .B(\u_div/PartRem[16][3] ), .Y(
        \u_div/u_add_PartRem_2_15/n3 ) );
  OR2X1 U353 ( .A(\u_div/PartRem[15][5] ), .B(\u_div/u_add_PartRem_2_14/n2 ), 
        .Y(\u_div/CryTmp[14][6] ) );
  XNOR2X1 U354 ( .A(\u_div/PartRem[15][3] ), .B(\u_div/PartRem[15][2] ), .Y(
        \u_div/SumTmp[14][3] ) );
  XNOR2X1 U355 ( .A(\u_div/PartRem[14][3] ), .B(\u_div/PartRem[14][2] ), .Y(
        \u_div/SumTmp[13][3] ) );
  OR2X1 U356 ( .A(\u_div/PartRem[14][2] ), .B(\u_div/PartRem[14][3] ), .Y(
        \u_div/u_add_PartRem_2_13/n3 ) );
  OR2X1 U357 ( .A(\u_div/PartRem[13][5] ), .B(\u_div/u_add_PartRem_2_12/n2 ), 
        .Y(\u_div/CryTmp[12][6] ) );
  XNOR2X1 U358 ( .A(\u_div/PartRem[13][3] ), .B(\u_div/PartRem[13][2] ), .Y(
        \u_div/SumTmp[12][3] ) );
  XNOR2X1 U359 ( .A(\u_div/PartRem[12][3] ), .B(\u_div/PartRem[12][2] ), .Y(
        \u_div/SumTmp[11][3] ) );
  XNOR2X1 U360 ( .A(\u_div/PartRem[11][3] ), .B(\u_div/PartRem[11][2] ), .Y(
        \u_div/SumTmp[10][3] ) );
  OR2X1 U361 ( .A(\u_div/PartRem[11][2] ), .B(\u_div/PartRem[11][3] ), .Y(
        \u_div/u_add_PartRem_2_10/n3 ) );
  XNOR2X1 U362 ( .A(\u_div/PartRem[10][3] ), .B(\u_div/PartRem[10][2] ), .Y(
        \u_div/SumTmp[9][3] ) );
  XNOR2X1 U363 ( .A(\u_div/PartRem[9][3] ), .B(\u_div/PartRem[9][2] ), .Y(
        \u_div/SumTmp[8][3] ) );
  OR2X1 U364 ( .A(\u_div/PartRem[9][2] ), .B(\u_div/PartRem[9][3] ), .Y(
        \u_div/u_add_PartRem_2_8/n3 ) );
  OR2X1 U365 ( .A(\u_div/PartRem[8][5] ), .B(\u_div/u_add_PartRem_2_7/n2 ), 
        .Y(\u_div/CryTmp[7][6] ) );
  XNOR2X1 U366 ( .A(\u_div/PartRem[8][3] ), .B(\u_div/PartRem[8][2] ), .Y(
        \u_div/SumTmp[7][3] ) );
  XNOR2X1 U367 ( .A(\u_div/PartRem[7][3] ), .B(\u_div/PartRem[7][2] ), .Y(
        \u_div/SumTmp[6][3] ) );
  XNOR2X1 U368 ( .A(\u_div/PartRem[6][3] ), .B(\u_div/PartRem[6][2] ), .Y(
        \u_div/SumTmp[5][3] ) );
  OR2X1 U369 ( .A(\u_div/PartRem[6][2] ), .B(\u_div/PartRem[6][3] ), .Y(
        \u_div/u_add_PartRem_2_5/n3 ) );
  XNOR2X1 U370 ( .A(\u_div/PartRem[5][3] ), .B(\u_div/PartRem[5][2] ), .Y(
        \u_div/SumTmp[4][3] ) );
  XNOR2X1 U371 ( .A(\u_div/PartRem[4][3] ), .B(\u_div/PartRem[4][2] ), .Y(
        \u_div/SumTmp[3][3] ) );
  OR2X1 U372 ( .A(\u_div/PartRem[4][2] ), .B(\u_div/PartRem[4][3] ), .Y(
        \u_div/u_add_PartRem_2_3/n3 ) );
  XNOR2X1 U373 ( .A(\u_div/PartRem[3][3] ), .B(\u_div/PartRem[3][2] ), .Y(
        \u_div/SumTmp[2][3] ) );
  XNOR2X1 U374 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/PartRem[2][2] ), .Y(
        \u_div/SumTmp[1][3] ) );
  OR2X1 U375 ( .A(\u_div/PartRem[2][2] ), .B(\u_div/PartRem[2][3] ), .Y(
        \u_div/u_add_PartRem_2_1/n3 ) );
  XNOR2X1 U376 ( .A(\u_div/PartRem[63][0] ), .B(\u_div/PartRem[62][0] ), .Y(
        \u_div/SumTmp[59][3] ) );
  XOR2X1 U377 ( .A(\u_div/CryTmp[8][6] ), .B(n7), .Y(\u_div/QInv[8] ) );
  XOR2X1 U378 ( .A(\u_div/CryTmp[7][6] ), .B(n8), .Y(\u_div/QInv[7] ) );
  XOR2X1 U379 ( .A(\u_div/CryTmp[59][6] ), .B(n7), .Y(\u_div/QInv[59] ) );
  XOR2X1 U380 ( .A(\u_div/CryTmp[58][6] ), .B(n9), .Y(\u_div/QInv[58] ) );
  XOR2X1 U381 ( .A(\u_div/CryTmp[57][6] ), .B(n8), .Y(\u_div/QInv[57] ) );
  XOR2X1 U382 ( .A(\u_div/CryTmp[56][6] ), .B(n7), .Y(\u_div/QInv[56] ) );
  XOR2X1 U383 ( .A(\u_div/CryTmp[55][6] ), .B(n9), .Y(\u_div/QInv[55] ) );
  XOR2X1 U384 ( .A(\u_div/CryTmp[51][6] ), .B(n8), .Y(\u_div/QInv[51] ) );
  XOR2X1 U385 ( .A(\u_div/CryTmp[50][6] ), .B(n7), .Y(\u_div/QInv[50] ) );
  XOR2X1 U386 ( .A(\u_div/CryTmp[49][6] ), .B(n8), .Y(\u_div/QInv[49] ) );
  XOR2X1 U387 ( .A(\u_div/CryTmp[48][6] ), .B(n7), .Y(\u_div/QInv[48] ) );
  XOR2X1 U388 ( .A(\u_div/CryTmp[47][6] ), .B(n9), .Y(\u_div/QInv[47] ) );
  XOR2X1 U389 ( .A(\u_div/CryTmp[43][6] ), .B(n8), .Y(\u_div/QInv[43] ) );
  XOR2X1 U390 ( .A(\u_div/CryTmp[42][6] ), .B(n7), .Y(\u_div/QInv[42] ) );
  XOR2X1 U391 ( .A(\u_div/CryTmp[41][6] ), .B(n9), .Y(\u_div/QInv[41] ) );
  XOR2X1 U392 ( .A(\u_div/CryTmp[40][6] ), .B(n8), .Y(\u_div/QInv[40] ) );
  XOR2X1 U393 ( .A(\u_div/CryTmp[3][6] ), .B(n7), .Y(\u_div/QInv[3] ) );
  XOR2X1 U394 ( .A(\u_div/CryTmp[39][6] ), .B(n9), .Y(\u_div/QInv[39] ) );
  XOR2X1 U395 ( .A(\u_div/CryTmp[38][6] ), .B(n8), .Y(\u_div/QInv[38] ) );
  XOR2X1 U396 ( .A(\u_div/CryTmp[37][6] ), .B(n7), .Y(\u_div/QInv[37] ) );
  XOR2X1 U397 ( .A(\u_div/CryTmp[33][6] ), .B(n8), .Y(\u_div/QInv[33] ) );
  XOR2X1 U398 ( .A(\u_div/CryTmp[32][6] ), .B(n7), .Y(\u_div/QInv[32] ) );
  XOR2X1 U399 ( .A(\u_div/CryTmp[31][6] ), .B(n9), .Y(\u_div/QInv[31] ) );
  XOR2X1 U400 ( .A(\u_div/CryTmp[30][6] ), .B(n8), .Y(\u_div/QInv[30] ) );
  XOR2X1 U401 ( .A(\u_div/CryTmp[2][6] ), .B(n7), .Y(\u_div/QInv[2] ) );
  XOR2X1 U402 ( .A(\u_div/CryTmp[29][6] ), .B(n9), .Y(\u_div/QInv[29] ) );
  XOR2X1 U403 ( .A(\u_div/CryTmp[28][6] ), .B(n8), .Y(\u_div/QInv[28] ) );
  XOR2X1 U404 ( .A(\u_div/CryTmp[27][6] ), .B(n7), .Y(\u_div/QInv[27] ) );
  XOR2X1 U405 ( .A(\u_div/CryTmp[23][6] ), .B(n9), .Y(\u_div/QInv[23] ) );
  XOR2X1 U406 ( .A(\u_div/CryTmp[22][6] ), .B(n8), .Y(\u_div/QInv[22] ) );
  XOR2X1 U407 ( .A(\u_div/CryTmp[20][6] ), .B(n9), .Y(\u_div/QInv[20] ) );
  XOR2X1 U408 ( .A(\u_div/CryTmp[1][6] ), .B(n8), .Y(\u_div/QInv[1] ) );
  XOR2X1 U409 ( .A(\u_div/CryTmp[18][6] ), .B(n9), .Y(\u_div/QInv[18] ) );
  XOR2X1 U410 ( .A(\u_div/CryTmp[17][6] ), .B(n8), .Y(\u_div/QInv[17] ) );
  XOR2X1 U411 ( .A(\u_div/CryTmp[13][6] ), .B(n8), .Y(\u_div/QInv[13] ) );
  XOR2X1 U412 ( .A(\u_div/CryTmp[12][6] ), .B(n9), .Y(\u_div/QInv[12] ) );
  XOR2X1 U413 ( .A(\u_div/CryTmp[11][6] ), .B(n8), .Y(\u_div/QInv[11] ) );
  XOR2X1 U414 ( .A(\u_div/CryTmp[10][6] ), .B(n9), .Y(\u_div/QInv[10] ) );
endmodule


module GSIM_DW01_inc_9 ( A, SUM );
  input [63:0] A;
  output [63:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58;

  NOR3BX1 U2 ( .AN(A[59]), .B(n1), .C(n17), .Y(n15) );
  NAND3X1 U3 ( .A(A[56]), .B(n19), .C(A[57]), .Y(n17) );
  NOR3BX1 U4 ( .AN(A[19]), .B(n11), .C(n57), .Y(n55) );
  NOR3BX1 U5 ( .AN(A[51]), .B(n3), .C(n25), .Y(n23) );
  NAND3X1 U6 ( .A(A[48]), .B(n27), .C(A[49]), .Y(n25) );
  NOR3BX1 U7 ( .AN(A[43]), .B(n5), .C(n33), .Y(n31) );
  NAND3X1 U8 ( .A(A[40]), .B(n35), .C(A[41]), .Y(n33) );
  NOR3BX1 U9 ( .AN(A[35]), .B(n7), .C(n41), .Y(n39) );
  NAND3X1 U10 ( .A(A[32]), .B(n43), .C(A[33]), .Y(n41) );
  NOR3BX1 U11 ( .AN(A[27]), .B(n9), .C(n49), .Y(n47) );
  NAND3X1 U12 ( .A(A[24]), .B(n51), .C(A[25]), .Y(n49) );
  NOR3BX1 U13 ( .AN(A[47]), .B(n4), .C(n29), .Y(n27) );
  NOR3BX1 U14 ( .AN(A[39]), .B(n6), .C(n37), .Y(n35) );
  NOR3BX1 U15 ( .AN(A[31]), .B(n8), .C(n45), .Y(n43) );
  NOR3BX1 U16 ( .AN(A[23]), .B(n10), .C(n53), .Y(n51) );
  NOR3BX1 U17 ( .AN(A[55]), .B(n2), .C(n21), .Y(n19) );
  NAND3XL U18 ( .A(A[60]), .B(n15), .C(A[61]), .Y(n14) );
  NAND3XL U19 ( .A(A[52]), .B(n23), .C(A[53]), .Y(n21) );
  NAND3XL U20 ( .A(A[44]), .B(n31), .C(A[45]), .Y(n29) );
  NAND3XL U21 ( .A(A[36]), .B(n39), .C(A[37]), .Y(n37) );
  NAND3XL U22 ( .A(A[28]), .B(n47), .C(A[29]), .Y(n45) );
  NAND3XL U23 ( .A(A[20]), .B(n55), .C(A[21]), .Y(n53) );
  NAND2XL U24 ( .A(A[56]), .B(n19), .Y(n20) );
  NAND2XL U25 ( .A(A[52]), .B(n23), .Y(n24) );
  NAND2XL U26 ( .A(A[48]), .B(n27), .Y(n28) );
  NAND2XL U27 ( .A(A[44]), .B(n31), .Y(n32) );
  NAND2XL U28 ( .A(A[40]), .B(n35), .Y(n36) );
  NAND2XL U29 ( .A(A[36]), .B(n39), .Y(n40) );
  NAND2XL U30 ( .A(A[32]), .B(n43), .Y(n44) );
  NAND2XL U31 ( .A(A[28]), .B(n47), .Y(n48) );
  NAND2XL U32 ( .A(A[24]), .B(n51), .Y(n52) );
  NAND2XL U33 ( .A(A[20]), .B(n55), .Y(n56) );
  XOR2XL U34 ( .A(A[60]), .B(n15), .Y(SUM[60]) );
  NAND2XL U35 ( .A(A[60]), .B(n15), .Y(n16) );
  CLKINVX1 U36 ( .A(A[16]), .Y(SUM[16]) );
  CLKINVX1 U37 ( .A(A[18]), .Y(n11) );
  CLKINVX1 U38 ( .A(A[22]), .Y(n10) );
  CLKINVX1 U39 ( .A(A[26]), .Y(n9) );
  CLKINVX1 U40 ( .A(A[30]), .Y(n8) );
  CLKINVX1 U41 ( .A(A[34]), .Y(n7) );
  CLKINVX1 U42 ( .A(A[38]), .Y(n6) );
  CLKINVX1 U43 ( .A(A[42]), .Y(n5) );
  CLKINVX1 U44 ( .A(A[46]), .Y(n4) );
  CLKINVX1 U45 ( .A(A[50]), .Y(n3) );
  CLKINVX1 U46 ( .A(A[54]), .Y(n2) );
  CLKINVX1 U47 ( .A(A[58]), .Y(n1) );
  XOR2X1 U48 ( .A(A[63]), .B(n13), .Y(SUM[63]) );
  NOR2BX1 U49 ( .AN(A[62]), .B(n14), .Y(n13) );
  XNOR2X1 U50 ( .A(A[62]), .B(n14), .Y(SUM[62]) );
  XNOR2X1 U51 ( .A(A[61]), .B(n16), .Y(SUM[61]) );
  XOR2X1 U52 ( .A(A[59]), .B(n18), .Y(SUM[59]) );
  NOR2X1 U53 ( .A(n17), .B(n1), .Y(n18) );
  XOR2X1 U54 ( .A(n1), .B(n17), .Y(SUM[58]) );
  XNOR2X1 U55 ( .A(A[57]), .B(n20), .Y(SUM[57]) );
  XOR2X1 U56 ( .A(A[56]), .B(n19), .Y(SUM[56]) );
  XOR2X1 U57 ( .A(A[55]), .B(n22), .Y(SUM[55]) );
  NOR2X1 U58 ( .A(n21), .B(n2), .Y(n22) );
  XOR2X1 U59 ( .A(n2), .B(n21), .Y(SUM[54]) );
  XNOR2X1 U60 ( .A(A[53]), .B(n24), .Y(SUM[53]) );
  XOR2X1 U61 ( .A(A[52]), .B(n23), .Y(SUM[52]) );
  XOR2X1 U62 ( .A(A[51]), .B(n26), .Y(SUM[51]) );
  NOR2X1 U63 ( .A(n25), .B(n3), .Y(n26) );
  XOR2X1 U64 ( .A(n3), .B(n25), .Y(SUM[50]) );
  XNOR2X1 U65 ( .A(A[49]), .B(n28), .Y(SUM[49]) );
  XOR2X1 U66 ( .A(A[48]), .B(n27), .Y(SUM[48]) );
  XOR2X1 U67 ( .A(A[47]), .B(n30), .Y(SUM[47]) );
  NOR2X1 U68 ( .A(n29), .B(n4), .Y(n30) );
  XOR2X1 U69 ( .A(n4), .B(n29), .Y(SUM[46]) );
  XNOR2X1 U70 ( .A(A[45]), .B(n32), .Y(SUM[45]) );
  XOR2X1 U71 ( .A(A[44]), .B(n31), .Y(SUM[44]) );
  XOR2X1 U72 ( .A(A[43]), .B(n34), .Y(SUM[43]) );
  NOR2X1 U73 ( .A(n33), .B(n5), .Y(n34) );
  XOR2X1 U74 ( .A(n5), .B(n33), .Y(SUM[42]) );
  XNOR2X1 U75 ( .A(A[41]), .B(n36), .Y(SUM[41]) );
  XOR2X1 U76 ( .A(A[40]), .B(n35), .Y(SUM[40]) );
  XOR2X1 U77 ( .A(A[39]), .B(n38), .Y(SUM[39]) );
  NOR2X1 U78 ( .A(n37), .B(n6), .Y(n38) );
  XOR2X1 U79 ( .A(n6), .B(n37), .Y(SUM[38]) );
  XNOR2X1 U80 ( .A(A[37]), .B(n40), .Y(SUM[37]) );
  XOR2X1 U81 ( .A(A[36]), .B(n39), .Y(SUM[36]) );
  XOR2X1 U82 ( .A(A[35]), .B(n42), .Y(SUM[35]) );
  NOR2X1 U83 ( .A(n41), .B(n7), .Y(n42) );
  XOR2X1 U84 ( .A(n7), .B(n41), .Y(SUM[34]) );
  XNOR2X1 U85 ( .A(A[33]), .B(n44), .Y(SUM[33]) );
  XOR2X1 U86 ( .A(A[32]), .B(n43), .Y(SUM[32]) );
  XOR2X1 U87 ( .A(A[31]), .B(n46), .Y(SUM[31]) );
  NOR2X1 U88 ( .A(n45), .B(n8), .Y(n46) );
  XOR2X1 U89 ( .A(n8), .B(n45), .Y(SUM[30]) );
  XNOR2X1 U90 ( .A(A[29]), .B(n48), .Y(SUM[29]) );
  XOR2X1 U91 ( .A(A[28]), .B(n47), .Y(SUM[28]) );
  XOR2X1 U92 ( .A(A[27]), .B(n50), .Y(SUM[27]) );
  NOR2X1 U93 ( .A(n49), .B(n9), .Y(n50) );
  XOR2X1 U94 ( .A(n9), .B(n49), .Y(SUM[26]) );
  XNOR2X1 U95 ( .A(A[25]), .B(n52), .Y(SUM[25]) );
  XOR2X1 U96 ( .A(A[24]), .B(n51), .Y(SUM[24]) );
  XOR2X1 U97 ( .A(A[23]), .B(n54), .Y(SUM[23]) );
  NOR2X1 U98 ( .A(n53), .B(n10), .Y(n54) );
  XOR2X1 U99 ( .A(n10), .B(n53), .Y(SUM[22]) );
  XNOR2X1 U100 ( .A(A[21]), .B(n56), .Y(SUM[21]) );
  XOR2X1 U101 ( .A(A[20]), .B(n55), .Y(SUM[20]) );
  XOR2X1 U102 ( .A(A[19]), .B(n58), .Y(SUM[19]) );
  NOR2X1 U103 ( .A(n57), .B(n11), .Y(n58) );
  XOR2X1 U104 ( .A(n11), .B(n57), .Y(SUM[18]) );
  NAND2X1 U105 ( .A(A[17]), .B(A[16]), .Y(n57) );
  XOR2X1 U106 ( .A(A[17]), .B(A[16]), .Y(SUM[17]) );
endmodule


module GSIM_DW01_absval_7 ( A, ABSVAL );
  input [63:0] A;
  output [63:0] ABSVAL;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51;
  wire   [63:0] AMUX1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  GSIM_DW01_inc_9 NEG ( .A({n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
        n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .SUM({AMUX1[63:16], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15}) );
  AND2X2 U1 ( .A(AMUX1[63]), .B(n3), .Y(ABSVAL[63]) );
  CLKINVX1 U2 ( .A(A[63]), .Y(n4) );
  INVX3 U3 ( .A(n4), .Y(n3) );
  INVX3 U4 ( .A(n4), .Y(n2) );
  INVX3 U5 ( .A(n4), .Y(n1) );
  CLKINVX1 U6 ( .A(A[16]), .Y(n51) );
  CLKINVX1 U7 ( .A(A[17]), .Y(n50) );
  CLKINVX1 U8 ( .A(A[18]), .Y(n49) );
  CLKINVX1 U9 ( .A(A[19]), .Y(n48) );
  CLKINVX1 U10 ( .A(A[20]), .Y(n47) );
  CLKINVX1 U11 ( .A(A[21]), .Y(n46) );
  CLKINVX1 U12 ( .A(A[22]), .Y(n45) );
  CLKINVX1 U13 ( .A(A[23]), .Y(n44) );
  CLKINVX1 U14 ( .A(A[24]), .Y(n43) );
  CLKINVX1 U15 ( .A(A[25]), .Y(n42) );
  CLKINVX1 U16 ( .A(A[26]), .Y(n41) );
  CLKINVX1 U17 ( .A(A[27]), .Y(n40) );
  CLKINVX1 U18 ( .A(A[28]), .Y(n39) );
  CLKINVX1 U19 ( .A(A[29]), .Y(n38) );
  CLKINVX1 U20 ( .A(A[30]), .Y(n37) );
  CLKINVX1 U21 ( .A(A[31]), .Y(n36) );
  CLKINVX1 U22 ( .A(A[32]), .Y(n35) );
  CLKINVX1 U23 ( .A(A[33]), .Y(n34) );
  CLKINVX1 U24 ( .A(A[34]), .Y(n33) );
  CLKINVX1 U25 ( .A(A[35]), .Y(n32) );
  CLKINVX1 U26 ( .A(A[36]), .Y(n31) );
  CLKINVX1 U27 ( .A(A[37]), .Y(n30) );
  CLKINVX1 U28 ( .A(A[38]), .Y(n29) );
  CLKINVX1 U29 ( .A(A[39]), .Y(n28) );
  CLKINVX1 U30 ( .A(A[40]), .Y(n27) );
  CLKINVX1 U31 ( .A(A[41]), .Y(n26) );
  CLKINVX1 U32 ( .A(A[42]), .Y(n25) );
  CLKINVX1 U33 ( .A(A[43]), .Y(n24) );
  CLKINVX1 U34 ( .A(A[44]), .Y(n23) );
  CLKINVX1 U35 ( .A(A[45]), .Y(n22) );
  CLKINVX1 U36 ( .A(A[46]), .Y(n21) );
  CLKINVX1 U37 ( .A(A[47]), .Y(n20) );
  CLKINVX1 U38 ( .A(A[48]), .Y(n19) );
  CLKINVX1 U39 ( .A(A[49]), .Y(n18) );
  CLKINVX1 U40 ( .A(A[50]), .Y(n17) );
  CLKINVX1 U41 ( .A(A[51]), .Y(n16) );
  CLKINVX1 U42 ( .A(A[52]), .Y(n15) );
  CLKINVX1 U43 ( .A(A[53]), .Y(n14) );
  CLKINVX1 U44 ( .A(A[54]), .Y(n13) );
  CLKINVX1 U45 ( .A(A[55]), .Y(n12) );
  CLKINVX1 U46 ( .A(A[56]), .Y(n11) );
  CLKINVX1 U47 ( .A(A[57]), .Y(n10) );
  CLKINVX1 U48 ( .A(A[58]), .Y(n9) );
  CLKINVX1 U49 ( .A(A[59]), .Y(n8) );
  CLKINVX1 U50 ( .A(A[60]), .Y(n7) );
  CLKINVX1 U51 ( .A(A[61]), .Y(n6) );
  CLKINVX1 U52 ( .A(A[62]), .Y(n5) );
  CLKMX2X2 U54 ( .A(A[62]), .B(AMUX1[62]), .S0(n3), .Y(ABSVAL[62]) );
  CLKMX2X2 U55 ( .A(A[61]), .B(AMUX1[61]), .S0(n3), .Y(ABSVAL[61]) );
  CLKMX2X2 U56 ( .A(A[60]), .B(AMUX1[60]), .S0(n3), .Y(ABSVAL[60]) );
  CLKMX2X2 U57 ( .A(A[59]), .B(AMUX1[59]), .S0(n3), .Y(ABSVAL[59]) );
  CLKMX2X2 U58 ( .A(A[58]), .B(AMUX1[58]), .S0(n3), .Y(ABSVAL[58]) );
  CLKMX2X2 U59 ( .A(A[57]), .B(AMUX1[57]), .S0(n3), .Y(ABSVAL[57]) );
  CLKMX2X2 U60 ( .A(A[56]), .B(AMUX1[56]), .S0(n3), .Y(ABSVAL[56]) );
  CLKMX2X2 U61 ( .A(A[55]), .B(AMUX1[55]), .S0(n3), .Y(ABSVAL[55]) );
  CLKMX2X2 U62 ( .A(A[54]), .B(AMUX1[54]), .S0(n2), .Y(ABSVAL[54]) );
  CLKMX2X2 U63 ( .A(A[53]), .B(AMUX1[53]), .S0(n2), .Y(ABSVAL[53]) );
  CLKMX2X2 U64 ( .A(A[52]), .B(AMUX1[52]), .S0(n2), .Y(ABSVAL[52]) );
  CLKMX2X2 U65 ( .A(A[51]), .B(AMUX1[51]), .S0(n2), .Y(ABSVAL[51]) );
  CLKMX2X2 U66 ( .A(A[50]), .B(AMUX1[50]), .S0(n2), .Y(ABSVAL[50]) );
  CLKMX2X2 U67 ( .A(A[49]), .B(AMUX1[49]), .S0(n2), .Y(ABSVAL[49]) );
  CLKMX2X2 U68 ( .A(A[48]), .B(AMUX1[48]), .S0(n2), .Y(ABSVAL[48]) );
  CLKMX2X2 U69 ( .A(A[47]), .B(AMUX1[47]), .S0(n2), .Y(ABSVAL[47]) );
  CLKMX2X2 U70 ( .A(A[46]), .B(AMUX1[46]), .S0(n2), .Y(ABSVAL[46]) );
  CLKMX2X2 U71 ( .A(A[45]), .B(AMUX1[45]), .S0(n2), .Y(ABSVAL[45]) );
  CLKMX2X2 U72 ( .A(A[44]), .B(AMUX1[44]), .S0(n2), .Y(ABSVAL[44]) );
  CLKMX2X2 U73 ( .A(A[43]), .B(AMUX1[43]), .S0(n2), .Y(ABSVAL[43]) );
  CLKMX2X2 U74 ( .A(A[42]), .B(AMUX1[42]), .S0(n2), .Y(ABSVAL[42]) );
  CLKMX2X2 U75 ( .A(A[41]), .B(AMUX1[41]), .S0(n1), .Y(ABSVAL[41]) );
  CLKMX2X2 U76 ( .A(A[40]), .B(AMUX1[40]), .S0(n1), .Y(ABSVAL[40]) );
  CLKMX2X2 U77 ( .A(A[39]), .B(AMUX1[39]), .S0(n1), .Y(ABSVAL[39]) );
  CLKMX2X2 U78 ( .A(A[38]), .B(AMUX1[38]), .S0(n1), .Y(ABSVAL[38]) );
  CLKMX2X2 U79 ( .A(A[37]), .B(AMUX1[37]), .S0(n1), .Y(ABSVAL[37]) );
  CLKMX2X2 U80 ( .A(A[36]), .B(AMUX1[36]), .S0(n1), .Y(ABSVAL[36]) );
  CLKMX2X2 U81 ( .A(A[35]), .B(AMUX1[35]), .S0(n1), .Y(ABSVAL[35]) );
  CLKMX2X2 U82 ( .A(A[34]), .B(AMUX1[34]), .S0(n1), .Y(ABSVAL[34]) );
  CLKMX2X2 U83 ( .A(A[33]), .B(AMUX1[33]), .S0(n1), .Y(ABSVAL[33]) );
  CLKMX2X2 U84 ( .A(A[32]), .B(AMUX1[32]), .S0(n1), .Y(ABSVAL[32]) );
  CLKMX2X2 U85 ( .A(A[31]), .B(AMUX1[31]), .S0(n1), .Y(ABSVAL[31]) );
  CLKMX2X2 U86 ( .A(A[30]), .B(AMUX1[30]), .S0(n1), .Y(ABSVAL[30]) );
  CLKMX2X2 U87 ( .A(A[29]), .B(AMUX1[29]), .S0(n1), .Y(ABSVAL[29]) );
  CLKMX2X2 U88 ( .A(A[28]), .B(AMUX1[28]), .S0(n1), .Y(ABSVAL[28]) );
  CLKMX2X2 U89 ( .A(A[27]), .B(AMUX1[27]), .S0(n1), .Y(ABSVAL[27]) );
  CLKMX2X2 U90 ( .A(A[26]), .B(AMUX1[26]), .S0(n1), .Y(ABSVAL[26]) );
  CLKMX2X2 U91 ( .A(A[25]), .B(AMUX1[25]), .S0(n1), .Y(ABSVAL[25]) );
  CLKMX2X2 U92 ( .A(A[24]), .B(AMUX1[24]), .S0(n2), .Y(ABSVAL[24]) );
  CLKMX2X2 U93 ( .A(A[23]), .B(AMUX1[23]), .S0(n2), .Y(ABSVAL[23]) );
  CLKMX2X2 U94 ( .A(A[22]), .B(AMUX1[22]), .S0(n2), .Y(ABSVAL[22]) );
  CLKMX2X2 U95 ( .A(A[21]), .B(AMUX1[21]), .S0(n2), .Y(ABSVAL[21]) );
  CLKMX2X2 U96 ( .A(A[20]), .B(AMUX1[20]), .S0(n3), .Y(ABSVAL[20]) );
  CLKMX2X2 U97 ( .A(A[19]), .B(AMUX1[19]), .S0(n3), .Y(ABSVAL[19]) );
  CLKMX2X2 U98 ( .A(A[18]), .B(AMUX1[18]), .S0(n3), .Y(ABSVAL[18]) );
  CLKMX2X2 U99 ( .A(A[17]), .B(AMUX1[17]), .S0(n3), .Y(ABSVAL[17]) );
  CLKMX2X2 U100 ( .A(A[16]), .B(AMUX1[16]), .S0(n3), .Y(ABSVAL[16]) );
endmodule


module GSIM_DW_inc_7 ( carry_in, a, carry_out, sum );
  input [63:0] a;
  output [63:0] sum;
  input carry_in;
  output carry_out;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63;

  ADDHXL U7 ( .A(a[59]), .B(n5), .CO(n4), .S(sum[59]) );
  ADDHXL U8 ( .A(a[58]), .B(n6), .CO(n5), .S(sum[58]) );
  ADDHXL U9 ( .A(a[57]), .B(n7), .CO(n6), .S(sum[57]) );
  ADDHXL U10 ( .A(a[56]), .B(n8), .CO(n7), .S(sum[56]) );
  ADDHXL U11 ( .A(a[55]), .B(n9), .CO(n8), .S(sum[55]) );
  ADDHXL U12 ( .A(a[54]), .B(n10), .CO(n9), .S(sum[54]) );
  ADDHXL U13 ( .A(a[53]), .B(n11), .CO(n10), .S(sum[53]) );
  ADDHXL U14 ( .A(a[52]), .B(n12), .CO(n11), .S(sum[52]) );
  ADDHXL U15 ( .A(a[51]), .B(n13), .CO(n12), .S(sum[51]) );
  ADDHXL U16 ( .A(a[50]), .B(n14), .CO(n13), .S(sum[50]) );
  ADDHXL U17 ( .A(a[49]), .B(n15), .CO(n14), .S(sum[49]) );
  ADDHXL U18 ( .A(a[48]), .B(n16), .CO(n15), .S(sum[48]) );
  ADDHXL U19 ( .A(a[47]), .B(n17), .CO(n16), .S(sum[47]) );
  ADDHXL U20 ( .A(a[46]), .B(n18), .CO(n17), .S(sum[46]) );
  ADDHXL U21 ( .A(a[45]), .B(n19), .CO(n18), .S(sum[45]) );
  ADDHXL U22 ( .A(a[44]), .B(n20), .CO(n19), .S(sum[44]) );
  ADDHXL U23 ( .A(a[43]), .B(n21), .CO(n20), .S(sum[43]) );
  ADDHXL U24 ( .A(a[42]), .B(n22), .CO(n21), .S(sum[42]) );
  ADDHXL U25 ( .A(a[41]), .B(n23), .CO(n22), .S(sum[41]) );
  ADDHXL U26 ( .A(a[40]), .B(n24), .CO(n23), .S(sum[40]) );
  ADDHXL U27 ( .A(a[39]), .B(n25), .CO(n24), .S(sum[39]) );
  ADDHXL U28 ( .A(a[38]), .B(n26), .CO(n25), .S(sum[38]) );
  ADDHXL U29 ( .A(a[37]), .B(n27), .CO(n26), .S(sum[37]) );
  ADDHXL U30 ( .A(a[36]), .B(n28), .CO(n27), .S(sum[36]) );
  ADDHXL U31 ( .A(a[35]), .B(n29), .CO(n28), .S(sum[35]) );
  ADDHXL U32 ( .A(a[34]), .B(n30), .CO(n29), .S(sum[34]) );
  ADDHXL U33 ( .A(a[33]), .B(n31), .CO(n30), .S(sum[33]) );
  ADDHXL U34 ( .A(a[32]), .B(n32), .CO(n31), .S(sum[32]) );
  ADDHXL U35 ( .A(a[31]), .B(n33), .CO(n32), .S(sum[31]) );
  ADDHXL U36 ( .A(a[30]), .B(n34), .CO(n33), .S(sum[30]) );
  ADDHXL U37 ( .A(a[29]), .B(n35), .CO(n34), .S(sum[29]) );
  ADDHXL U38 ( .A(a[28]), .B(n36), .CO(n35), .S(sum[28]) );
  ADDHXL U39 ( .A(a[27]), .B(n37), .CO(n36), .S(sum[27]) );
  ADDHXL U40 ( .A(a[26]), .B(n38), .CO(n37), .S(sum[26]) );
  ADDHXL U41 ( .A(a[25]), .B(n39), .CO(n38), .S(sum[25]) );
  ADDHXL U42 ( .A(a[24]), .B(n40), .CO(n39), .S(sum[24]) );
  ADDHXL U43 ( .A(a[23]), .B(n41), .CO(n40), .S(sum[23]) );
  ADDHXL U44 ( .A(a[22]), .B(n42), .CO(n41), .S(sum[22]) );
  ADDHXL U45 ( .A(a[21]), .B(n43), .CO(n42), .S(sum[21]) );
  ADDHXL U46 ( .A(a[20]), .B(n44), .CO(n43), .S(sum[20]) );
  ADDHXL U47 ( .A(a[19]), .B(n45), .CO(n44), .S(sum[19]) );
  ADDHXL U48 ( .A(a[18]), .B(n46), .CO(n45), .S(sum[18]) );
  ADDHXL U49 ( .A(a[17]), .B(n47), .CO(n46), .S(sum[17]) );
  ADDHXL U50 ( .A(a[16]), .B(n48), .CO(n47), .S(sum[16]) );
  ADDHXL U51 ( .A(a[15]), .B(n49), .CO(n48), .S(sum[15]) );
  ADDHXL U52 ( .A(a[14]), .B(n50), .CO(n49), .S(sum[14]) );
  ADDHXL U53 ( .A(a[13]), .B(n51), .CO(n50), .S(sum[13]) );
  ADDHXL U54 ( .A(a[12]), .B(n52), .CO(n51), .S(sum[12]) );
  ADDHXL U55 ( .A(a[11]), .B(n53), .CO(n52), .S(sum[11]) );
  ADDHXL U56 ( .A(a[10]), .B(n54), .CO(n53), .S(sum[10]) );
  ADDHXL U57 ( .A(a[9]), .B(n55), .CO(n54), .S(sum[9]) );
  ADDHXL U58 ( .A(a[8]), .B(n56), .CO(n55), .S(sum[8]) );
  ADDHXL U59 ( .A(a[7]), .B(n57), .CO(n56), .S(sum[7]) );
  ADDHXL U60 ( .A(a[6]), .B(n58), .CO(n57), .S(sum[6]) );
  ADDHXL U61 ( .A(a[5]), .B(n59), .CO(n58), .S(sum[5]) );
  ADDHXL U62 ( .A(a[4]), .B(n60), .CO(n59), .S(sum[4]) );
  ADDHXL U63 ( .A(a[3]), .B(n61), .CO(n60), .S(sum[3]) );
  ADDHXL U64 ( .A(a[2]), .B(n62), .CO(n61), .S(sum[2]) );
  ADDHXL U65 ( .A(a[1]), .B(n63), .CO(n62), .S(sum[1]) );
  ADDHXL U66 ( .A(carry_in), .B(a[0]), .CO(n63), .S(sum[0]) );
  NOR2BX1 U70 ( .AN(a[61]), .B(n4), .Y(sum[63]) );
  XOR2X1 U71 ( .A(a[61]), .B(n4), .Y(sum[60]) );
endmodule


module GSIM_DW_div_tc_7 ( a, b, quotient, remainder, divide_by_0 );
  input [63:0] a;
  input [5:0] b;
  output [63:0] quotient;
  output [5:0] remainder;
  output divide_by_0;
  wire   \u_div/QInv[63] , \u_div/QInv[59] , \u_div/QInv[58] ,
         \u_div/QInv[57] , \u_div/QInv[56] , \u_div/QInv[55] ,
         \u_div/QInv[54] , \u_div/QInv[53] , \u_div/QInv[52] ,
         \u_div/QInv[51] , \u_div/QInv[50] , \u_div/QInv[49] ,
         \u_div/QInv[48] , \u_div/QInv[47] , \u_div/QInv[46] ,
         \u_div/QInv[45] , \u_div/QInv[44] , \u_div/QInv[43] ,
         \u_div/QInv[42] , \u_div/QInv[41] , \u_div/QInv[40] ,
         \u_div/QInv[39] , \u_div/QInv[38] , \u_div/QInv[37] ,
         \u_div/QInv[36] , \u_div/QInv[35] , \u_div/QInv[34] ,
         \u_div/QInv[33] , \u_div/QInv[32] , \u_div/QInv[31] ,
         \u_div/QInv[30] , \u_div/QInv[29] , \u_div/QInv[28] ,
         \u_div/QInv[27] , \u_div/QInv[26] , \u_div/QInv[25] ,
         \u_div/QInv[24] , \u_div/QInv[23] , \u_div/QInv[22] ,
         \u_div/QInv[21] , \u_div/QInv[20] , \u_div/QInv[19] ,
         \u_div/QInv[18] , \u_div/QInv[17] , \u_div/QInv[16] ,
         \u_div/QInv[15] , \u_div/QInv[14] , \u_div/QInv[13] ,
         \u_div/QInv[12] , \u_div/QInv[11] , \u_div/QInv[10] , \u_div/QInv[9] ,
         \u_div/QInv[8] , \u_div/QInv[7] , \u_div/QInv[6] , \u_div/QInv[5] ,
         \u_div/QInv[4] , \u_div/QInv[3] , \u_div/QInv[2] , \u_div/QInv[1] ,
         \u_div/QInv[0] , \u_div/SumTmp[1][3] , \u_div/SumTmp[1][4] ,
         \u_div/SumTmp[2][3] , \u_div/SumTmp[2][4] , \u_div/SumTmp[3][3] ,
         \u_div/SumTmp[3][4] , \u_div/SumTmp[4][3] , \u_div/SumTmp[4][4] ,
         \u_div/SumTmp[5][3] , \u_div/SumTmp[5][4] , \u_div/SumTmp[6][3] ,
         \u_div/SumTmp[6][4] , \u_div/SumTmp[7][3] , \u_div/SumTmp[7][4] ,
         \u_div/SumTmp[8][3] , \u_div/SumTmp[8][4] , \u_div/SumTmp[9][3] ,
         \u_div/SumTmp[9][4] , \u_div/SumTmp[10][3] , \u_div/SumTmp[10][4] ,
         \u_div/SumTmp[11][3] , \u_div/SumTmp[11][4] , \u_div/SumTmp[12][3] ,
         \u_div/SumTmp[12][4] , \u_div/SumTmp[13][3] , \u_div/SumTmp[13][4] ,
         \u_div/SumTmp[14][2] , \u_div/SumTmp[14][3] , \u_div/SumTmp[14][4] ,
         \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] , \u_div/SumTmp[15][3] ,
         \u_div/SumTmp[15][4] , \u_div/SumTmp[16][1] , \u_div/SumTmp[16][2] ,
         \u_div/SumTmp[16][3] , \u_div/SumTmp[16][4] , \u_div/SumTmp[17][1] ,
         \u_div/SumTmp[17][2] , \u_div/SumTmp[17][3] , \u_div/SumTmp[17][4] ,
         \u_div/SumTmp[18][1] , \u_div/SumTmp[18][2] , \u_div/SumTmp[18][3] ,
         \u_div/SumTmp[18][4] , \u_div/SumTmp[19][1] , \u_div/SumTmp[19][2] ,
         \u_div/SumTmp[19][3] , \u_div/SumTmp[19][4] , \u_div/SumTmp[20][1] ,
         \u_div/SumTmp[20][2] , \u_div/SumTmp[20][3] , \u_div/SumTmp[20][4] ,
         \u_div/SumTmp[21][1] , \u_div/SumTmp[21][2] , \u_div/SumTmp[21][3] ,
         \u_div/SumTmp[21][4] , \u_div/SumTmp[22][1] , \u_div/SumTmp[22][2] ,
         \u_div/SumTmp[22][3] , \u_div/SumTmp[22][4] , \u_div/SumTmp[23][1] ,
         \u_div/SumTmp[23][2] , \u_div/SumTmp[23][3] , \u_div/SumTmp[23][4] ,
         \u_div/SumTmp[24][1] , \u_div/SumTmp[24][2] , \u_div/SumTmp[24][3] ,
         \u_div/SumTmp[24][4] , \u_div/SumTmp[25][1] , \u_div/SumTmp[25][2] ,
         \u_div/SumTmp[25][3] , \u_div/SumTmp[25][4] , \u_div/SumTmp[26][1] ,
         \u_div/SumTmp[26][2] , \u_div/SumTmp[26][3] , \u_div/SumTmp[26][4] ,
         \u_div/SumTmp[27][1] , \u_div/SumTmp[27][2] , \u_div/SumTmp[27][3] ,
         \u_div/SumTmp[27][4] , \u_div/SumTmp[28][1] , \u_div/SumTmp[28][2] ,
         \u_div/SumTmp[28][3] , \u_div/SumTmp[28][4] , \u_div/SumTmp[29][1] ,
         \u_div/SumTmp[29][2] , \u_div/SumTmp[29][3] , \u_div/SumTmp[29][4] ,
         \u_div/SumTmp[30][1] , \u_div/SumTmp[30][2] , \u_div/SumTmp[30][3] ,
         \u_div/SumTmp[30][4] , \u_div/SumTmp[31][1] , \u_div/SumTmp[31][2] ,
         \u_div/SumTmp[31][3] , \u_div/SumTmp[31][4] , \u_div/SumTmp[32][1] ,
         \u_div/SumTmp[32][2] , \u_div/SumTmp[32][3] , \u_div/SumTmp[32][4] ,
         \u_div/SumTmp[33][1] , \u_div/SumTmp[33][2] , \u_div/SumTmp[33][3] ,
         \u_div/SumTmp[33][4] , \u_div/SumTmp[34][1] , \u_div/SumTmp[34][2] ,
         \u_div/SumTmp[34][3] , \u_div/SumTmp[34][4] , \u_div/SumTmp[35][1] ,
         \u_div/SumTmp[35][2] , \u_div/SumTmp[35][3] , \u_div/SumTmp[35][4] ,
         \u_div/SumTmp[36][1] , \u_div/SumTmp[36][2] , \u_div/SumTmp[36][3] ,
         \u_div/SumTmp[36][4] , \u_div/SumTmp[37][1] , \u_div/SumTmp[37][2] ,
         \u_div/SumTmp[37][3] , \u_div/SumTmp[37][4] , \u_div/SumTmp[38][1] ,
         \u_div/SumTmp[38][2] , \u_div/SumTmp[38][3] , \u_div/SumTmp[38][4] ,
         \u_div/SumTmp[39][1] , \u_div/SumTmp[39][2] , \u_div/SumTmp[39][3] ,
         \u_div/SumTmp[39][4] , \u_div/SumTmp[40][1] , \u_div/SumTmp[40][2] ,
         \u_div/SumTmp[40][3] , \u_div/SumTmp[40][4] , \u_div/SumTmp[41][1] ,
         \u_div/SumTmp[41][2] , \u_div/SumTmp[41][3] , \u_div/SumTmp[41][4] ,
         \u_div/SumTmp[42][1] , \u_div/SumTmp[42][2] , \u_div/SumTmp[42][3] ,
         \u_div/SumTmp[42][4] , \u_div/SumTmp[43][1] , \u_div/SumTmp[43][2] ,
         \u_div/SumTmp[43][3] , \u_div/SumTmp[43][4] , \u_div/SumTmp[44][1] ,
         \u_div/SumTmp[44][2] , \u_div/SumTmp[44][3] , \u_div/SumTmp[44][4] ,
         \u_div/SumTmp[45][1] , \u_div/SumTmp[45][2] , \u_div/SumTmp[45][3] ,
         \u_div/SumTmp[45][4] , \u_div/SumTmp[46][1] , \u_div/SumTmp[46][2] ,
         \u_div/SumTmp[46][3] , \u_div/SumTmp[46][4] , \u_div/SumTmp[47][1] ,
         \u_div/SumTmp[47][2] , \u_div/SumTmp[47][3] , \u_div/SumTmp[47][4] ,
         \u_div/SumTmp[48][1] , \u_div/SumTmp[48][2] , \u_div/SumTmp[48][3] ,
         \u_div/SumTmp[48][4] , \u_div/SumTmp[49][1] , \u_div/SumTmp[49][2] ,
         \u_div/SumTmp[49][3] , \u_div/SumTmp[49][4] , \u_div/SumTmp[50][1] ,
         \u_div/SumTmp[50][2] , \u_div/SumTmp[50][3] , \u_div/SumTmp[50][4] ,
         \u_div/SumTmp[51][1] , \u_div/SumTmp[51][2] , \u_div/SumTmp[51][3] ,
         \u_div/SumTmp[51][4] , \u_div/SumTmp[52][1] , \u_div/SumTmp[52][2] ,
         \u_div/SumTmp[52][3] , \u_div/SumTmp[52][4] , \u_div/SumTmp[53][1] ,
         \u_div/SumTmp[53][2] , \u_div/SumTmp[53][3] , \u_div/SumTmp[53][4] ,
         \u_div/SumTmp[54][1] , \u_div/SumTmp[54][2] , \u_div/SumTmp[54][3] ,
         \u_div/SumTmp[54][4] , \u_div/SumTmp[55][1] , \u_div/SumTmp[55][2] ,
         \u_div/SumTmp[55][3] , \u_div/SumTmp[55][4] , \u_div/SumTmp[56][1] ,
         \u_div/SumTmp[56][2] , \u_div/SumTmp[56][3] , \u_div/SumTmp[56][4] ,
         \u_div/SumTmp[57][1] , \u_div/SumTmp[57][2] , \u_div/SumTmp[57][3] ,
         \u_div/SumTmp[57][4] , \u_div/SumTmp[58][1] , \u_div/SumTmp[58][2] ,
         \u_div/SumTmp[58][3] , \u_div/SumTmp[58][4] , \u_div/SumTmp[59][3] ,
         \u_div/SumTmp[59][4] , \u_div/CryTmp[0][6] , \u_div/CryTmp[1][6] ,
         \u_div/CryTmp[2][6] , \u_div/CryTmp[3][6] , \u_div/CryTmp[4][6] ,
         \u_div/CryTmp[5][6] , \u_div/CryTmp[6][6] , \u_div/CryTmp[7][6] ,
         \u_div/CryTmp[8][6] , \u_div/CryTmp[9][6] , \u_div/CryTmp[10][6] ,
         \u_div/CryTmp[11][6] , \u_div/CryTmp[12][6] , \u_div/CryTmp[13][6] ,
         \u_div/CryTmp[14][6] , \u_div/CryTmp[15][6] , \u_div/CryTmp[16][6] ,
         \u_div/CryTmp[17][6] , \u_div/CryTmp[18][6] , \u_div/CryTmp[19][6] ,
         \u_div/CryTmp[20][6] , \u_div/CryTmp[21][6] , \u_div/CryTmp[22][6] ,
         \u_div/CryTmp[23][6] , \u_div/CryTmp[24][6] , \u_div/CryTmp[25][6] ,
         \u_div/CryTmp[26][6] , \u_div/CryTmp[27][6] , \u_div/CryTmp[28][6] ,
         \u_div/CryTmp[29][6] , \u_div/CryTmp[30][6] , \u_div/CryTmp[31][6] ,
         \u_div/CryTmp[32][6] , \u_div/CryTmp[33][6] , \u_div/CryTmp[34][6] ,
         \u_div/CryTmp[35][6] , \u_div/CryTmp[36][6] , \u_div/CryTmp[37][6] ,
         \u_div/CryTmp[38][6] , \u_div/CryTmp[39][6] , \u_div/CryTmp[40][6] ,
         \u_div/CryTmp[41][6] , \u_div/CryTmp[42][6] , \u_div/CryTmp[43][6] ,
         \u_div/CryTmp[44][6] , \u_div/CryTmp[45][6] , \u_div/CryTmp[46][6] ,
         \u_div/CryTmp[47][6] , \u_div/CryTmp[48][6] , \u_div/CryTmp[49][6] ,
         \u_div/CryTmp[50][6] , \u_div/CryTmp[51][6] , \u_div/CryTmp[52][6] ,
         \u_div/CryTmp[53][6] , \u_div/CryTmp[54][6] , \u_div/CryTmp[55][6] ,
         \u_div/CryTmp[56][6] , \u_div/CryTmp[57][6] , \u_div/CryTmp[58][6] ,
         \u_div/CryTmp[59][6] , \u_div/PartRem[1][4] , \u_div/PartRem[1][5] ,
         \u_div/PartRem[2][4] , \u_div/PartRem[2][5] , \u_div/PartRem[3][4] ,
         \u_div/PartRem[3][5] , \u_div/PartRem[4][4] , \u_div/PartRem[4][5] ,
         \u_div/PartRem[5][4] , \u_div/PartRem[5][5] , \u_div/PartRem[6][4] ,
         \u_div/PartRem[6][5] , \u_div/PartRem[7][4] , \u_div/PartRem[7][5] ,
         \u_div/PartRem[8][4] , \u_div/PartRem[8][5] , \u_div/PartRem[9][4] ,
         \u_div/PartRem[9][5] , \u_div/PartRem[10][4] , \u_div/PartRem[10][5] ,
         \u_div/PartRem[11][4] , \u_div/PartRem[11][5] ,
         \u_div/PartRem[12][4] , \u_div/PartRem[12][5] ,
         \u_div/PartRem[13][4] , \u_div/PartRem[13][5] ,
         \u_div/PartRem[14][3] , \u_div/PartRem[14][4] ,
         \u_div/PartRem[14][5] , \u_div/PartRem[15][2] ,
         \u_div/PartRem[15][3] , \u_div/PartRem[15][4] ,
         \u_div/PartRem[15][5] , \u_div/PartRem[16][2] ,
         \u_div/PartRem[16][3] , \u_div/PartRem[16][4] ,
         \u_div/PartRem[16][5] , \u_div/PartRem[17][0] ,
         \u_div/PartRem[17][2] , \u_div/PartRem[17][3] ,
         \u_div/PartRem[17][4] , \u_div/PartRem[17][5] ,
         \u_div/PartRem[18][0] , \u_div/PartRem[18][2] ,
         \u_div/PartRem[18][3] , \u_div/PartRem[18][4] ,
         \u_div/PartRem[18][5] , \u_div/PartRem[19][0] ,
         \u_div/PartRem[19][2] , \u_div/PartRem[19][3] ,
         \u_div/PartRem[19][4] , \u_div/PartRem[19][5] ,
         \u_div/PartRem[20][0] , \u_div/PartRem[20][2] ,
         \u_div/PartRem[20][3] , \u_div/PartRem[20][4] ,
         \u_div/PartRem[20][5] , \u_div/PartRem[21][0] ,
         \u_div/PartRem[21][2] , \u_div/PartRem[21][3] ,
         \u_div/PartRem[21][4] , \u_div/PartRem[21][5] ,
         \u_div/PartRem[22][0] , \u_div/PartRem[22][2] ,
         \u_div/PartRem[22][3] , \u_div/PartRem[22][4] ,
         \u_div/PartRem[22][5] , \u_div/PartRem[23][0] ,
         \u_div/PartRem[23][2] , \u_div/PartRem[23][3] ,
         \u_div/PartRem[23][4] , \u_div/PartRem[23][5] ,
         \u_div/PartRem[24][0] , \u_div/PartRem[24][2] ,
         \u_div/PartRem[24][3] , \u_div/PartRem[24][4] ,
         \u_div/PartRem[24][5] , \u_div/PartRem[25][0] ,
         \u_div/PartRem[25][2] , \u_div/PartRem[25][3] ,
         \u_div/PartRem[25][4] , \u_div/PartRem[25][5] ,
         \u_div/PartRem[26][0] , \u_div/PartRem[26][2] ,
         \u_div/PartRem[26][3] , \u_div/PartRem[26][4] ,
         \u_div/PartRem[26][5] , \u_div/PartRem[27][0] ,
         \u_div/PartRem[27][2] , \u_div/PartRem[27][3] ,
         \u_div/PartRem[27][4] , \u_div/PartRem[27][5] ,
         \u_div/PartRem[28][0] , \u_div/PartRem[28][2] ,
         \u_div/PartRem[28][3] , \u_div/PartRem[28][4] ,
         \u_div/PartRem[28][5] , \u_div/PartRem[29][0] ,
         \u_div/PartRem[29][2] , \u_div/PartRem[29][3] ,
         \u_div/PartRem[29][4] , \u_div/PartRem[29][5] ,
         \u_div/PartRem[30][0] , \u_div/PartRem[30][2] ,
         \u_div/PartRem[30][3] , \u_div/PartRem[30][4] ,
         \u_div/PartRem[30][5] , \u_div/PartRem[31][0] ,
         \u_div/PartRem[31][2] , \u_div/PartRem[31][3] ,
         \u_div/PartRem[31][4] , \u_div/PartRem[31][5] ,
         \u_div/PartRem[32][0] , \u_div/PartRem[32][2] ,
         \u_div/PartRem[32][3] , \u_div/PartRem[32][4] ,
         \u_div/PartRem[32][5] , \u_div/PartRem[33][0] ,
         \u_div/PartRem[33][2] , \u_div/PartRem[33][3] ,
         \u_div/PartRem[33][4] , \u_div/PartRem[33][5] ,
         \u_div/PartRem[34][0] , \u_div/PartRem[34][2] ,
         \u_div/PartRem[34][3] , \u_div/PartRem[34][4] ,
         \u_div/PartRem[34][5] , \u_div/PartRem[35][0] ,
         \u_div/PartRem[35][2] , \u_div/PartRem[35][3] ,
         \u_div/PartRem[35][4] , \u_div/PartRem[35][5] ,
         \u_div/PartRem[36][0] , \u_div/PartRem[36][2] ,
         \u_div/PartRem[36][3] , \u_div/PartRem[36][4] ,
         \u_div/PartRem[36][5] , \u_div/PartRem[37][0] ,
         \u_div/PartRem[37][2] , \u_div/PartRem[37][3] ,
         \u_div/PartRem[37][4] , \u_div/PartRem[37][5] ,
         \u_div/PartRem[38][0] , \u_div/PartRem[38][2] ,
         \u_div/PartRem[38][3] , \u_div/PartRem[38][4] ,
         \u_div/PartRem[38][5] , \u_div/PartRem[39][0] ,
         \u_div/PartRem[39][2] , \u_div/PartRem[39][3] ,
         \u_div/PartRem[39][4] , \u_div/PartRem[39][5] ,
         \u_div/PartRem[40][0] , \u_div/PartRem[40][2] ,
         \u_div/PartRem[40][3] , \u_div/PartRem[40][4] ,
         \u_div/PartRem[40][5] , \u_div/PartRem[41][0] ,
         \u_div/PartRem[41][2] , \u_div/PartRem[41][3] ,
         \u_div/PartRem[41][4] , \u_div/PartRem[41][5] ,
         \u_div/PartRem[42][0] , \u_div/PartRem[42][2] ,
         \u_div/PartRem[42][3] , \u_div/PartRem[42][4] ,
         \u_div/PartRem[42][5] , \u_div/PartRem[43][0] ,
         \u_div/PartRem[43][2] , \u_div/PartRem[43][3] ,
         \u_div/PartRem[43][4] , \u_div/PartRem[43][5] ,
         \u_div/PartRem[44][0] , \u_div/PartRem[44][2] ,
         \u_div/PartRem[44][3] , \u_div/PartRem[44][4] ,
         \u_div/PartRem[44][5] , \u_div/PartRem[45][0] ,
         \u_div/PartRem[45][2] , \u_div/PartRem[45][3] ,
         \u_div/PartRem[45][4] , \u_div/PartRem[45][5] ,
         \u_div/PartRem[46][0] , \u_div/PartRem[46][2] ,
         \u_div/PartRem[46][3] , \u_div/PartRem[46][4] ,
         \u_div/PartRem[46][5] , \u_div/PartRem[47][0] ,
         \u_div/PartRem[47][2] , \u_div/PartRem[47][3] ,
         \u_div/PartRem[47][4] , \u_div/PartRem[47][5] ,
         \u_div/PartRem[48][0] , \u_div/PartRem[48][2] ,
         \u_div/PartRem[48][3] , \u_div/PartRem[48][4] ,
         \u_div/PartRem[48][5] , \u_div/PartRem[49][0] ,
         \u_div/PartRem[49][2] , \u_div/PartRem[49][3] ,
         \u_div/PartRem[49][4] , \u_div/PartRem[49][5] ,
         \u_div/PartRem[50][0] , \u_div/PartRem[50][2] ,
         \u_div/PartRem[50][3] , \u_div/PartRem[50][4] ,
         \u_div/PartRem[50][5] , \u_div/PartRem[51][0] ,
         \u_div/PartRem[51][2] , \u_div/PartRem[51][3] ,
         \u_div/PartRem[51][4] , \u_div/PartRem[51][5] ,
         \u_div/PartRem[52][0] , \u_div/PartRem[52][2] ,
         \u_div/PartRem[52][3] , \u_div/PartRem[52][4] ,
         \u_div/PartRem[52][5] , \u_div/PartRem[53][0] ,
         \u_div/PartRem[53][2] , \u_div/PartRem[53][3] ,
         \u_div/PartRem[53][4] , \u_div/PartRem[53][5] ,
         \u_div/PartRem[54][0] , \u_div/PartRem[54][2] ,
         \u_div/PartRem[54][3] , \u_div/PartRem[54][4] ,
         \u_div/PartRem[54][5] , \u_div/PartRem[55][0] ,
         \u_div/PartRem[55][2] , \u_div/PartRem[55][3] ,
         \u_div/PartRem[55][4] , \u_div/PartRem[55][5] ,
         \u_div/PartRem[56][0] , \u_div/PartRem[56][2] ,
         \u_div/PartRem[56][3] , \u_div/PartRem[56][4] ,
         \u_div/PartRem[56][5] , \u_div/PartRem[57][0] ,
         \u_div/PartRem[57][2] , \u_div/PartRem[57][3] ,
         \u_div/PartRem[57][4] , \u_div/PartRem[57][5] ,
         \u_div/PartRem[58][0] , \u_div/PartRem[58][2] ,
         \u_div/PartRem[58][3] , \u_div/PartRem[58][4] ,
         \u_div/PartRem[58][5] , \u_div/PartRem[59][0] ,
         \u_div/PartRem[59][2] , \u_div/PartRem[59][3] ,
         \u_div/PartRem[59][4] , \u_div/PartRem[59][5] ,
         \u_div/PartRem[60][0] , \u_div/PartRem[61][0] ,
         \u_div/PartRem[62][0] , \u_div/PartRem[63][0] ,
         \u_div/PartRem[64][0] , \u_div/u_add_PartRem_2_1/n2 ,
         \u_div/u_add_PartRem_2_2/n2 , \u_div/u_add_PartRem_2_3/n2 ,
         \u_div/u_add_PartRem_2_4/n2 , \u_div/u_add_PartRem_2_5/n2 ,
         \u_div/u_add_PartRem_2_6/n2 , \u_div/u_add_PartRem_2_7/n2 ,
         \u_div/u_add_PartRem_2_8/n2 , \u_div/u_add_PartRem_2_9/n2 ,
         \u_div/u_add_PartRem_2_10/n2 , \u_div/u_add_PartRem_2_11/n2 ,
         \u_div/u_add_PartRem_2_12/n2 , \u_div/u_add_PartRem_2_13/n2 ,
         \u_div/u_add_PartRem_2_14/n3 , \u_div/u_add_PartRem_2_14/n2 ,
         \u_div/u_add_PartRem_2_15/n3 , \u_div/u_add_PartRem_2_15/n2 ,
         \u_div/u_add_PartRem_2_16/n3 , \u_div/u_add_PartRem_2_16/n2 ,
         \u_div/u_add_PartRem_2_17/n3 , \u_div/u_add_PartRem_2_17/n2 ,
         \u_div/u_add_PartRem_2_18/n3 , \u_div/u_add_PartRem_2_18/n2 ,
         \u_div/u_add_PartRem_2_19/n3 , \u_div/u_add_PartRem_2_19/n2 ,
         \u_div/u_add_PartRem_2_20/n3 , \u_div/u_add_PartRem_2_20/n2 ,
         \u_div/u_add_PartRem_2_21/n3 , \u_div/u_add_PartRem_2_21/n2 ,
         \u_div/u_add_PartRem_2_22/n3 , \u_div/u_add_PartRem_2_22/n2 ,
         \u_div/u_add_PartRem_2_23/n3 , \u_div/u_add_PartRem_2_23/n2 ,
         \u_div/u_add_PartRem_2_24/n3 , \u_div/u_add_PartRem_2_24/n2 ,
         \u_div/u_add_PartRem_2_25/n3 , \u_div/u_add_PartRem_2_25/n2 ,
         \u_div/u_add_PartRem_2_26/n3 , \u_div/u_add_PartRem_2_26/n2 ,
         \u_div/u_add_PartRem_2_27/n3 , \u_div/u_add_PartRem_2_27/n2 ,
         \u_div/u_add_PartRem_2_28/n3 , \u_div/u_add_PartRem_2_28/n2 ,
         \u_div/u_add_PartRem_2_29/n3 , \u_div/u_add_PartRem_2_29/n2 ,
         \u_div/u_add_PartRem_2_30/n3 , \u_div/u_add_PartRem_2_30/n2 ,
         \u_div/u_add_PartRem_2_31/n3 , \u_div/u_add_PartRem_2_31/n2 ,
         \u_div/u_add_PartRem_2_32/n3 , \u_div/u_add_PartRem_2_32/n2 ,
         \u_div/u_add_PartRem_2_33/n3 , \u_div/u_add_PartRem_2_33/n2 ,
         \u_div/u_add_PartRem_2_34/n3 , \u_div/u_add_PartRem_2_34/n2 ,
         \u_div/u_add_PartRem_2_35/n3 , \u_div/u_add_PartRem_2_35/n2 ,
         \u_div/u_add_PartRem_2_36/n3 , \u_div/u_add_PartRem_2_36/n2 ,
         \u_div/u_add_PartRem_2_37/n3 , \u_div/u_add_PartRem_2_37/n2 ,
         \u_div/u_add_PartRem_2_38/n3 , \u_div/u_add_PartRem_2_38/n2 ,
         \u_div/u_add_PartRem_2_39/n3 , \u_div/u_add_PartRem_2_39/n2 ,
         \u_div/u_add_PartRem_2_40/n3 , \u_div/u_add_PartRem_2_40/n2 ,
         \u_div/u_add_PartRem_2_41/n3 , \u_div/u_add_PartRem_2_41/n2 ,
         \u_div/u_add_PartRem_2_42/n3 , \u_div/u_add_PartRem_2_42/n2 ,
         \u_div/u_add_PartRem_2_43/n3 , \u_div/u_add_PartRem_2_43/n2 ,
         \u_div/u_add_PartRem_2_44/n3 , \u_div/u_add_PartRem_2_44/n2 ,
         \u_div/u_add_PartRem_2_45/n3 , \u_div/u_add_PartRem_2_45/n2 ,
         \u_div/u_add_PartRem_2_46/n3 , \u_div/u_add_PartRem_2_46/n2 ,
         \u_div/u_add_PartRem_2_47/n3 , \u_div/u_add_PartRem_2_47/n2 ,
         \u_div/u_add_PartRem_2_48/n3 , \u_div/u_add_PartRem_2_48/n2 ,
         \u_div/u_add_PartRem_2_49/n3 , \u_div/u_add_PartRem_2_49/n2 ,
         \u_div/u_add_PartRem_2_50/n3 , \u_div/u_add_PartRem_2_50/n2 ,
         \u_div/u_add_PartRem_2_51/n3 , \u_div/u_add_PartRem_2_51/n2 ,
         \u_div/u_add_PartRem_2_52/n3 , \u_div/u_add_PartRem_2_52/n2 ,
         \u_div/u_add_PartRem_2_53/n3 , \u_div/u_add_PartRem_2_53/n2 ,
         \u_div/u_add_PartRem_2_54/n3 , \u_div/u_add_PartRem_2_54/n2 ,
         \u_div/u_add_PartRem_2_55/n3 , \u_div/u_add_PartRem_2_55/n2 ,
         \u_div/u_add_PartRem_2_56/n3 , \u_div/u_add_PartRem_2_56/n2 ,
         \u_div/u_add_PartRem_2_57/n3 , \u_div/u_add_PartRem_2_57/n2 ,
         \u_div/u_add_PartRem_2_58/n3 , \u_div/u_add_PartRem_2_58/n2 , n1, n2,
         n3, n4, n5, n6;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17;
  assign \u_div/QInv[63]  = a[63];

  GSIM_DW01_absval_7 \u_div/u_absval_AAbs  ( .A({n2, a[62:16], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .ABSVAL({\u_div/PartRem[64][0] , \u_div/PartRem[63][0] , 
        \u_div/PartRem[62][0] , \u_div/PartRem[61][0] , \u_div/PartRem[60][0] , 
        \u_div/PartRem[59][0] , \u_div/PartRem[58][0] , \u_div/PartRem[57][0] , 
        \u_div/PartRem[56][0] , \u_div/PartRem[55][0] , \u_div/PartRem[54][0] , 
        \u_div/PartRem[53][0] , \u_div/PartRem[52][0] , \u_div/PartRem[51][0] , 
        \u_div/PartRem[50][0] , \u_div/PartRem[49][0] , \u_div/PartRem[48][0] , 
        \u_div/PartRem[47][0] , \u_div/PartRem[46][0] , \u_div/PartRem[45][0] , 
        \u_div/PartRem[44][0] , \u_div/PartRem[43][0] , \u_div/PartRem[42][0] , 
        \u_div/PartRem[41][0] , \u_div/PartRem[40][0] , \u_div/PartRem[39][0] , 
        \u_div/PartRem[38][0] , \u_div/PartRem[37][0] , \u_div/PartRem[36][0] , 
        \u_div/PartRem[35][0] , \u_div/PartRem[34][0] , \u_div/PartRem[33][0] , 
        \u_div/PartRem[32][0] , \u_div/PartRem[31][0] , \u_div/PartRem[30][0] , 
        \u_div/PartRem[29][0] , \u_div/PartRem[28][0] , \u_div/PartRem[27][0] , 
        \u_div/PartRem[26][0] , \u_div/PartRem[25][0] , \u_div/PartRem[24][0] , 
        \u_div/PartRem[23][0] , \u_div/PartRem[22][0] , \u_div/PartRem[21][0] , 
        \u_div/PartRem[20][0] , \u_div/PartRem[19][0] , \u_div/PartRem[18][0] , 
        \u_div/PartRem[17][0] , SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15}) );
  GSIM_DW_inc_7 \u_div/u_inc_QInc  ( .carry_in(n3), .a({n2, n2, 
        \u_div/QInv[63] , n2, \u_div/QInv[59] , \u_div/QInv[58] , 
        \u_div/QInv[57] , \u_div/QInv[56] , \u_div/QInv[55] , \u_div/QInv[54] , 
        \u_div/QInv[53] , \u_div/QInv[52] , \u_div/QInv[51] , \u_div/QInv[50] , 
        \u_div/QInv[49] , \u_div/QInv[48] , \u_div/QInv[47] , \u_div/QInv[46] , 
        \u_div/QInv[45] , \u_div/QInv[44] , \u_div/QInv[43] , \u_div/QInv[42] , 
        \u_div/QInv[41] , \u_div/QInv[40] , \u_div/QInv[39] , \u_div/QInv[38] , 
        \u_div/QInv[37] , \u_div/QInv[36] , \u_div/QInv[35] , \u_div/QInv[34] , 
        \u_div/QInv[33] , \u_div/QInv[32] , \u_div/QInv[31] , \u_div/QInv[30] , 
        \u_div/QInv[29] , \u_div/QInv[28] , \u_div/QInv[27] , \u_div/QInv[26] , 
        \u_div/QInv[25] , \u_div/QInv[24] , \u_div/QInv[23] , \u_div/QInv[22] , 
        \u_div/QInv[21] , \u_div/QInv[20] , \u_div/QInv[19] , \u_div/QInv[18] , 
        \u_div/QInv[17] , \u_div/QInv[16] , \u_div/QInv[15] , \u_div/QInv[14] , 
        \u_div/QInv[13] , \u_div/QInv[12] , \u_div/QInv[11] , \u_div/QInv[10] , 
        \u_div/QInv[9] , \u_div/QInv[8] , \u_div/QInv[7] , \u_div/QInv[6] , 
        \u_div/QInv[5] , \u_div/QInv[4] , \u_div/QInv[3] , \u_div/QInv[2] , 
        \u_div/QInv[1] , \u_div/QInv[0] }), .sum({quotient[63], 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, quotient[60:0]})
         );
  ADDHXL \u_div/u_add_PartRem_2_1/U3  ( .A(\u_div/PartRem[2][4] ), .B(
        \u_div/CryTmp[2][6] ), .CO(\u_div/u_add_PartRem_2_1/n2 ), .S(
        \u_div/SumTmp[1][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_2/U3  ( .A(\u_div/PartRem[3][4] ), .B(
        \u_div/CryTmp[3][6] ), .CO(\u_div/u_add_PartRem_2_2/n2 ), .S(
        \u_div/SumTmp[2][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_3/U3  ( .A(\u_div/PartRem[4][4] ), .B(
        \u_div/CryTmp[4][6] ), .CO(\u_div/u_add_PartRem_2_3/n2 ), .S(
        \u_div/SumTmp[3][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_4/U3  ( .A(\u_div/PartRem[5][4] ), .B(
        \u_div/CryTmp[5][6] ), .CO(\u_div/u_add_PartRem_2_4/n2 ), .S(
        \u_div/SumTmp[4][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_5/U3  ( .A(\u_div/PartRem[6][4] ), .B(
        \u_div/CryTmp[6][6] ), .CO(\u_div/u_add_PartRem_2_5/n2 ), .S(
        \u_div/SumTmp[5][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_6/U3  ( .A(\u_div/PartRem[7][4] ), .B(
        \u_div/CryTmp[7][6] ), .CO(\u_div/u_add_PartRem_2_6/n2 ), .S(
        \u_div/SumTmp[6][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_7/U3  ( .A(\u_div/PartRem[8][4] ), .B(
        \u_div/CryTmp[8][6] ), .CO(\u_div/u_add_PartRem_2_7/n2 ), .S(
        \u_div/SumTmp[7][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_8/U3  ( .A(\u_div/PartRem[9][4] ), .B(
        \u_div/CryTmp[9][6] ), .CO(\u_div/u_add_PartRem_2_8/n2 ), .S(
        \u_div/SumTmp[8][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_9/U3  ( .A(\u_div/PartRem[10][4] ), .B(
        \u_div/CryTmp[10][6] ), .CO(\u_div/u_add_PartRem_2_9/n2 ), .S(
        \u_div/SumTmp[9][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_10/U3  ( .A(\u_div/PartRem[11][4] ), .B(
        \u_div/CryTmp[11][6] ), .CO(\u_div/u_add_PartRem_2_10/n2 ), .S(
        \u_div/SumTmp[10][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_11/U3  ( .A(\u_div/PartRem[12][4] ), .B(
        \u_div/CryTmp[12][6] ), .CO(\u_div/u_add_PartRem_2_11/n2 ), .S(
        \u_div/SumTmp[11][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_12/U3  ( .A(\u_div/PartRem[13][4] ), .B(
        \u_div/CryTmp[13][6] ), .CO(\u_div/u_add_PartRem_2_12/n2 ), .S(
        \u_div/SumTmp[12][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_13/U3  ( .A(\u_div/PartRem[14][4] ), .B(
        \u_div/PartRem[14][3] ), .CO(\u_div/u_add_PartRem_2_13/n2 ), .S(
        \u_div/SumTmp[13][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_14/U3  ( .A(\u_div/PartRem[15][4] ), .B(
        \u_div/u_add_PartRem_2_14/n3 ), .CO(\u_div/u_add_PartRem_2_14/n2 ), 
        .S(\u_div/SumTmp[14][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_15/U3  ( .A(\u_div/PartRem[16][4] ), .B(
        \u_div/u_add_PartRem_2_15/n3 ), .CO(\u_div/u_add_PartRem_2_15/n2 ), 
        .S(\u_div/SumTmp[15][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_16/U3  ( .A(\u_div/PartRem[17][4] ), .B(
        \u_div/u_add_PartRem_2_16/n3 ), .CO(\u_div/u_add_PartRem_2_16/n2 ), 
        .S(\u_div/SumTmp[16][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_17/U3  ( .A(\u_div/PartRem[18][4] ), .B(
        \u_div/u_add_PartRem_2_17/n3 ), .CO(\u_div/u_add_PartRem_2_17/n2 ), 
        .S(\u_div/SumTmp[17][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_18/U3  ( .A(\u_div/PartRem[19][4] ), .B(
        \u_div/u_add_PartRem_2_18/n3 ), .CO(\u_div/u_add_PartRem_2_18/n2 ), 
        .S(\u_div/SumTmp[18][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_19/U3  ( .A(\u_div/PartRem[20][4] ), .B(
        \u_div/u_add_PartRem_2_19/n3 ), .CO(\u_div/u_add_PartRem_2_19/n2 ), 
        .S(\u_div/SumTmp[19][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_20/U3  ( .A(\u_div/PartRem[21][4] ), .B(
        \u_div/u_add_PartRem_2_20/n3 ), .CO(\u_div/u_add_PartRem_2_20/n2 ), 
        .S(\u_div/SumTmp[20][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_21/U3  ( .A(\u_div/PartRem[22][4] ), .B(
        \u_div/u_add_PartRem_2_21/n3 ), .CO(\u_div/u_add_PartRem_2_21/n2 ), 
        .S(\u_div/SumTmp[21][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_22/U3  ( .A(\u_div/PartRem[23][4] ), .B(
        \u_div/u_add_PartRem_2_22/n3 ), .CO(\u_div/u_add_PartRem_2_22/n2 ), 
        .S(\u_div/SumTmp[22][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_23/U3  ( .A(\u_div/PartRem[24][4] ), .B(
        \u_div/u_add_PartRem_2_23/n3 ), .CO(\u_div/u_add_PartRem_2_23/n2 ), 
        .S(\u_div/SumTmp[23][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_24/U3  ( .A(\u_div/PartRem[25][4] ), .B(
        \u_div/u_add_PartRem_2_24/n3 ), .CO(\u_div/u_add_PartRem_2_24/n2 ), 
        .S(\u_div/SumTmp[24][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_25/U3  ( .A(\u_div/PartRem[26][4] ), .B(
        \u_div/u_add_PartRem_2_25/n3 ), .CO(\u_div/u_add_PartRem_2_25/n2 ), 
        .S(\u_div/SumTmp[25][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_26/U3  ( .A(\u_div/PartRem[27][4] ), .B(
        \u_div/u_add_PartRem_2_26/n3 ), .CO(\u_div/u_add_PartRem_2_26/n2 ), 
        .S(\u_div/SumTmp[26][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_27/U3  ( .A(\u_div/PartRem[28][4] ), .B(
        \u_div/u_add_PartRem_2_27/n3 ), .CO(\u_div/u_add_PartRem_2_27/n2 ), 
        .S(\u_div/SumTmp[27][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_28/U3  ( .A(\u_div/PartRem[29][4] ), .B(
        \u_div/u_add_PartRem_2_28/n3 ), .CO(\u_div/u_add_PartRem_2_28/n2 ), 
        .S(\u_div/SumTmp[28][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_29/U3  ( .A(\u_div/PartRem[30][4] ), .B(
        \u_div/u_add_PartRem_2_29/n3 ), .CO(\u_div/u_add_PartRem_2_29/n2 ), 
        .S(\u_div/SumTmp[29][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_30/U3  ( .A(\u_div/PartRem[31][4] ), .B(
        \u_div/u_add_PartRem_2_30/n3 ), .CO(\u_div/u_add_PartRem_2_30/n2 ), 
        .S(\u_div/SumTmp[30][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_31/U3  ( .A(\u_div/PartRem[32][4] ), .B(
        \u_div/u_add_PartRem_2_31/n3 ), .CO(\u_div/u_add_PartRem_2_31/n2 ), 
        .S(\u_div/SumTmp[31][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_32/U3  ( .A(\u_div/PartRem[33][4] ), .B(
        \u_div/u_add_PartRem_2_32/n3 ), .CO(\u_div/u_add_PartRem_2_32/n2 ), 
        .S(\u_div/SumTmp[32][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_33/U3  ( .A(\u_div/PartRem[34][4] ), .B(
        \u_div/u_add_PartRem_2_33/n3 ), .CO(\u_div/u_add_PartRem_2_33/n2 ), 
        .S(\u_div/SumTmp[33][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_34/U3  ( .A(\u_div/PartRem[35][4] ), .B(
        \u_div/u_add_PartRem_2_34/n3 ), .CO(\u_div/u_add_PartRem_2_34/n2 ), 
        .S(\u_div/SumTmp[34][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_35/U3  ( .A(\u_div/PartRem[36][4] ), .B(
        \u_div/u_add_PartRem_2_35/n3 ), .CO(\u_div/u_add_PartRem_2_35/n2 ), 
        .S(\u_div/SumTmp[35][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_36/U3  ( .A(\u_div/PartRem[37][4] ), .B(
        \u_div/u_add_PartRem_2_36/n3 ), .CO(\u_div/u_add_PartRem_2_36/n2 ), 
        .S(\u_div/SumTmp[36][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_37/U3  ( .A(\u_div/PartRem[38][4] ), .B(
        \u_div/u_add_PartRem_2_37/n3 ), .CO(\u_div/u_add_PartRem_2_37/n2 ), 
        .S(\u_div/SumTmp[37][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_38/U3  ( .A(\u_div/PartRem[39][4] ), .B(
        \u_div/u_add_PartRem_2_38/n3 ), .CO(\u_div/u_add_PartRem_2_38/n2 ), 
        .S(\u_div/SumTmp[38][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_39/U3  ( .A(\u_div/PartRem[40][4] ), .B(
        \u_div/u_add_PartRem_2_39/n3 ), .CO(\u_div/u_add_PartRem_2_39/n2 ), 
        .S(\u_div/SumTmp[39][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_40/U3  ( .A(\u_div/PartRem[41][4] ), .B(
        \u_div/u_add_PartRem_2_40/n3 ), .CO(\u_div/u_add_PartRem_2_40/n2 ), 
        .S(\u_div/SumTmp[40][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_41/U3  ( .A(\u_div/PartRem[42][4] ), .B(
        \u_div/u_add_PartRem_2_41/n3 ), .CO(\u_div/u_add_PartRem_2_41/n2 ), 
        .S(\u_div/SumTmp[41][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_42/U3  ( .A(\u_div/PartRem[43][4] ), .B(
        \u_div/u_add_PartRem_2_42/n3 ), .CO(\u_div/u_add_PartRem_2_42/n2 ), 
        .S(\u_div/SumTmp[42][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_43/U3  ( .A(\u_div/PartRem[44][4] ), .B(
        \u_div/u_add_PartRem_2_43/n3 ), .CO(\u_div/u_add_PartRem_2_43/n2 ), 
        .S(\u_div/SumTmp[43][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_44/U3  ( .A(\u_div/PartRem[45][4] ), .B(
        \u_div/u_add_PartRem_2_44/n3 ), .CO(\u_div/u_add_PartRem_2_44/n2 ), 
        .S(\u_div/SumTmp[44][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_45/U3  ( .A(\u_div/PartRem[46][4] ), .B(
        \u_div/u_add_PartRem_2_45/n3 ), .CO(\u_div/u_add_PartRem_2_45/n2 ), 
        .S(\u_div/SumTmp[45][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_46/U3  ( .A(\u_div/PartRem[47][4] ), .B(
        \u_div/u_add_PartRem_2_46/n3 ), .CO(\u_div/u_add_PartRem_2_46/n2 ), 
        .S(\u_div/SumTmp[46][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_47/U3  ( .A(\u_div/PartRem[48][4] ), .B(
        \u_div/u_add_PartRem_2_47/n3 ), .CO(\u_div/u_add_PartRem_2_47/n2 ), 
        .S(\u_div/SumTmp[47][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_48/U3  ( .A(\u_div/PartRem[49][4] ), .B(
        \u_div/u_add_PartRem_2_48/n3 ), .CO(\u_div/u_add_PartRem_2_48/n2 ), 
        .S(\u_div/SumTmp[48][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_49/U3  ( .A(\u_div/PartRem[50][4] ), .B(
        \u_div/u_add_PartRem_2_49/n3 ), .CO(\u_div/u_add_PartRem_2_49/n2 ), 
        .S(\u_div/SumTmp[49][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_50/U3  ( .A(\u_div/PartRem[51][4] ), .B(
        \u_div/u_add_PartRem_2_50/n3 ), .CO(\u_div/u_add_PartRem_2_50/n2 ), 
        .S(\u_div/SumTmp[50][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_51/U3  ( .A(\u_div/PartRem[52][4] ), .B(
        \u_div/u_add_PartRem_2_51/n3 ), .CO(\u_div/u_add_PartRem_2_51/n2 ), 
        .S(\u_div/SumTmp[51][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_52/U3  ( .A(\u_div/PartRem[53][4] ), .B(
        \u_div/u_add_PartRem_2_52/n3 ), .CO(\u_div/u_add_PartRem_2_52/n2 ), 
        .S(\u_div/SumTmp[52][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_53/U3  ( .A(\u_div/PartRem[54][4] ), .B(
        \u_div/u_add_PartRem_2_53/n3 ), .CO(\u_div/u_add_PartRem_2_53/n2 ), 
        .S(\u_div/SumTmp[53][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_54/U3  ( .A(\u_div/PartRem[55][4] ), .B(
        \u_div/u_add_PartRem_2_54/n3 ), .CO(\u_div/u_add_PartRem_2_54/n2 ), 
        .S(\u_div/SumTmp[54][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_55/U3  ( .A(\u_div/PartRem[56][4] ), .B(
        \u_div/u_add_PartRem_2_55/n3 ), .CO(\u_div/u_add_PartRem_2_55/n2 ), 
        .S(\u_div/SumTmp[55][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_56/U3  ( .A(\u_div/PartRem[57][4] ), .B(
        \u_div/u_add_PartRem_2_56/n3 ), .CO(\u_div/u_add_PartRem_2_56/n2 ), 
        .S(\u_div/SumTmp[56][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_57/U3  ( .A(\u_div/PartRem[58][4] ), .B(
        \u_div/u_add_PartRem_2_57/n3 ), .CO(\u_div/u_add_PartRem_2_57/n2 ), 
        .S(\u_div/SumTmp[57][4] ) );
  ADDHXL \u_div/u_add_PartRem_2_58/U3  ( .A(\u_div/PartRem[59][4] ), .B(
        \u_div/u_add_PartRem_2_58/n3 ), .CO(\u_div/u_add_PartRem_2_58/n2 ), 
        .S(\u_div/SumTmp[58][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_0  ( .A(\u_div/PartRem[17][0] ), .B(
        \u_div/PartRem[17][0] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/SumTmp[15][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_15_1  ( .A(\u_div/SumTmp[15][1] ), .B(
        \u_div/SumTmp[15][1] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_0  ( .A(\u_div/PartRem[18][0] ), .B(
        \u_div/PartRem[18][0] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/SumTmp[16][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_16_1  ( .A(\u_div/SumTmp[16][1] ), .B(
        \u_div/SumTmp[16][1] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_0  ( .A(\u_div/PartRem[19][0] ), .B(
        \u_div/PartRem[19][0] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/SumTmp[17][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_17_1  ( .A(\u_div/SumTmp[17][1] ), .B(
        \u_div/SumTmp[17][1] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_0  ( .A(\u_div/PartRem[20][0] ), .B(
        \u_div/PartRem[20][0] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/SumTmp[18][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_18_1  ( .A(\u_div/SumTmp[18][1] ), .B(
        \u_div/SumTmp[18][1] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_0  ( .A(\u_div/PartRem[21][0] ), .B(
        \u_div/PartRem[21][0] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/SumTmp[19][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_19_1  ( .A(\u_div/SumTmp[19][1] ), .B(
        \u_div/SumTmp[19][1] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_0  ( .A(\u_div/PartRem[22][0] ), .B(
        \u_div/PartRem[22][0] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/SumTmp[20][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_20_1  ( .A(\u_div/SumTmp[20][1] ), .B(
        \u_div/SumTmp[20][1] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_0  ( .A(\u_div/PartRem[23][0] ), .B(
        \u_div/PartRem[23][0] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/SumTmp[21][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_21_1  ( .A(\u_div/SumTmp[21][1] ), .B(
        \u_div/SumTmp[21][1] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_0  ( .A(\u_div/PartRem[24][0] ), .B(
        \u_div/PartRem[24][0] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/SumTmp[22][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_22_1  ( .A(\u_div/SumTmp[22][1] ), .B(
        \u_div/SumTmp[22][1] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_0  ( .A(\u_div/PartRem[25][0] ), .B(
        \u_div/PartRem[25][0] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/SumTmp[23][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_23_1  ( .A(\u_div/SumTmp[23][1] ), .B(
        \u_div/SumTmp[23][1] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_0  ( .A(\u_div/PartRem[26][0] ), .B(
        \u_div/PartRem[26][0] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/SumTmp[24][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_24_1  ( .A(\u_div/SumTmp[24][1] ), .B(
        \u_div/SumTmp[24][1] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_0  ( .A(\u_div/PartRem[27][0] ), .B(
        \u_div/PartRem[27][0] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/SumTmp[25][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_25_1  ( .A(\u_div/SumTmp[25][1] ), .B(
        \u_div/SumTmp[25][1] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_0  ( .A(\u_div/PartRem[28][0] ), .B(
        \u_div/PartRem[28][0] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/SumTmp[26][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_26_1  ( .A(\u_div/SumTmp[26][1] ), .B(
        \u_div/SumTmp[26][1] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_0  ( .A(\u_div/PartRem[29][0] ), .B(
        \u_div/PartRem[29][0] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/SumTmp[27][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_27_1  ( .A(\u_div/SumTmp[27][1] ), .B(
        \u_div/SumTmp[27][1] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_0  ( .A(\u_div/PartRem[30][0] ), .B(
        \u_div/PartRem[30][0] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/SumTmp[28][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_28_1  ( .A(\u_div/SumTmp[28][1] ), .B(
        \u_div/SumTmp[28][1] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_0  ( .A(\u_div/PartRem[31][0] ), .B(
        \u_div/PartRem[31][0] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/SumTmp[29][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_29_1  ( .A(\u_div/SumTmp[29][1] ), .B(
        \u_div/SumTmp[29][1] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_0  ( .A(\u_div/PartRem[32][0] ), .B(
        \u_div/PartRem[32][0] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/SumTmp[30][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_30_1  ( .A(\u_div/SumTmp[30][1] ), .B(
        \u_div/SumTmp[30][1] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_0  ( .A(\u_div/PartRem[33][0] ), .B(
        \u_div/PartRem[33][0] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/SumTmp[31][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_31_1  ( .A(\u_div/SumTmp[31][1] ), .B(
        \u_div/SumTmp[31][1] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_0  ( .A(\u_div/PartRem[34][0] ), .B(
        \u_div/PartRem[34][0] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/SumTmp[32][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_32_1  ( .A(\u_div/SumTmp[32][1] ), .B(
        \u_div/SumTmp[32][1] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_0  ( .A(\u_div/PartRem[35][0] ), .B(
        \u_div/PartRem[35][0] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/SumTmp[33][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_33_1  ( .A(\u_div/SumTmp[33][1] ), .B(
        \u_div/SumTmp[33][1] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_0  ( .A(\u_div/PartRem[36][0] ), .B(
        \u_div/PartRem[36][0] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/SumTmp[34][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_34_1  ( .A(\u_div/SumTmp[34][1] ), .B(
        \u_div/SumTmp[34][1] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_0  ( .A(\u_div/PartRem[37][0] ), .B(
        \u_div/PartRem[37][0] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/SumTmp[35][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_35_1  ( .A(\u_div/SumTmp[35][1] ), .B(
        \u_div/SumTmp[35][1] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_0  ( .A(\u_div/PartRem[38][0] ), .B(
        \u_div/PartRem[38][0] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/SumTmp[36][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_36_1  ( .A(\u_div/SumTmp[36][1] ), .B(
        \u_div/SumTmp[36][1] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_0  ( .A(\u_div/PartRem[39][0] ), .B(
        \u_div/PartRem[39][0] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/SumTmp[37][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_37_1  ( .A(\u_div/SumTmp[37][1] ), .B(
        \u_div/SumTmp[37][1] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_0  ( .A(\u_div/PartRem[40][0] ), .B(
        \u_div/PartRem[40][0] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/SumTmp[38][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_38_1  ( .A(\u_div/SumTmp[38][1] ), .B(
        \u_div/SumTmp[38][1] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_0  ( .A(\u_div/PartRem[41][0] ), .B(
        \u_div/PartRem[41][0] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/SumTmp[39][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_39_1  ( .A(\u_div/SumTmp[39][1] ), .B(
        \u_div/SumTmp[39][1] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_0  ( .A(\u_div/PartRem[42][0] ), .B(
        \u_div/PartRem[42][0] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/SumTmp[40][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_40_1  ( .A(\u_div/SumTmp[40][1] ), .B(
        \u_div/SumTmp[40][1] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_0  ( .A(\u_div/PartRem[43][0] ), .B(
        \u_div/PartRem[43][0] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/SumTmp[41][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_41_1  ( .A(\u_div/SumTmp[41][1] ), .B(
        \u_div/SumTmp[41][1] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_0  ( .A(\u_div/PartRem[44][0] ), .B(
        \u_div/PartRem[44][0] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/SumTmp[42][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_42_1  ( .A(\u_div/SumTmp[42][1] ), .B(
        \u_div/SumTmp[42][1] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_0  ( .A(\u_div/PartRem[45][0] ), .B(
        \u_div/PartRem[45][0] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/SumTmp[43][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_43_1  ( .A(\u_div/SumTmp[43][1] ), .B(
        \u_div/SumTmp[43][1] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_0  ( .A(\u_div/PartRem[46][0] ), .B(
        \u_div/PartRem[46][0] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/SumTmp[44][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_44_1  ( .A(\u_div/SumTmp[44][1] ), .B(
        \u_div/SumTmp[44][1] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_0  ( .A(\u_div/PartRem[47][0] ), .B(
        \u_div/PartRem[47][0] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/SumTmp[45][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_45_1  ( .A(\u_div/SumTmp[45][1] ), .B(
        \u_div/SumTmp[45][1] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_0  ( .A(\u_div/PartRem[48][0] ), .B(
        \u_div/PartRem[48][0] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/SumTmp[46][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_46_1  ( .A(\u_div/SumTmp[46][1] ), .B(
        \u_div/SumTmp[46][1] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_0  ( .A(\u_div/PartRem[49][0] ), .B(
        \u_div/PartRem[49][0] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/SumTmp[47][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_47_1  ( .A(\u_div/SumTmp[47][1] ), .B(
        \u_div/SumTmp[47][1] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_0  ( .A(\u_div/PartRem[50][0] ), .B(
        \u_div/PartRem[50][0] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/SumTmp[48][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_48_1  ( .A(\u_div/SumTmp[48][1] ), .B(
        \u_div/SumTmp[48][1] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_0  ( .A(\u_div/PartRem[51][0] ), .B(
        \u_div/PartRem[51][0] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/SumTmp[49][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_49_1  ( .A(\u_div/SumTmp[49][1] ), .B(
        \u_div/SumTmp[49][1] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_0  ( .A(\u_div/PartRem[52][0] ), .B(
        \u_div/PartRem[52][0] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/SumTmp[50][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_50_1  ( .A(\u_div/SumTmp[50][1] ), .B(
        \u_div/SumTmp[50][1] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_0  ( .A(\u_div/PartRem[53][0] ), .B(
        \u_div/PartRem[53][0] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/SumTmp[51][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_51_1  ( .A(\u_div/SumTmp[51][1] ), .B(
        \u_div/SumTmp[51][1] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_0  ( .A(\u_div/PartRem[54][0] ), .B(
        \u_div/PartRem[54][0] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/SumTmp[52][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_52_1  ( .A(\u_div/SumTmp[52][1] ), .B(
        \u_div/SumTmp[52][1] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_0  ( .A(\u_div/PartRem[55][0] ), .B(
        \u_div/PartRem[55][0] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/SumTmp[53][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_53_1  ( .A(\u_div/SumTmp[53][1] ), .B(
        \u_div/SumTmp[53][1] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_0  ( .A(\u_div/PartRem[56][0] ), .B(
        \u_div/PartRem[56][0] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/SumTmp[54][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_54_1  ( .A(\u_div/SumTmp[54][1] ), .B(
        \u_div/SumTmp[54][1] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_0  ( .A(\u_div/PartRem[57][0] ), .B(
        \u_div/PartRem[57][0] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/SumTmp[55][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_55_1  ( .A(\u_div/SumTmp[55][1] ), .B(
        \u_div/SumTmp[55][1] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_0  ( .A(\u_div/PartRem[58][0] ), .B(
        \u_div/PartRem[58][0] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/SumTmp[56][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_56_1  ( .A(\u_div/SumTmp[56][1] ), .B(
        \u_div/SumTmp[56][1] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_0  ( .A(\u_div/PartRem[59][0] ), .B(
        \u_div/PartRem[59][0] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/SumTmp[57][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_57_1  ( .A(\u_div/SumTmp[57][1] ), .B(
        \u_div/SumTmp[57][1] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][2] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_0  ( .A(\u_div/PartRem[60][0] ), .B(
        \u_div/PartRem[60][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/SumTmp[58][1] ) );
  MX2X1 \u_div/u_mx_PartRem_1_58_1  ( .A(\u_div/SumTmp[58][1] ), .B(
        \u_div/SumTmp[58][1] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][2] ) );
  MX2X1 \u_div/u_mx_PartRem_1_59_1  ( .A(\u_div/PartRem[61][0] ), .B(
        \u_div/PartRem[61][0] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_15_3  ( .A(\u_div/PartRem[16][3] ), .B(
        \u_div/SumTmp[15][3] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_16_3  ( .A(\u_div/PartRem[17][3] ), .B(
        \u_div/SumTmp[16][3] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_17_3  ( .A(\u_div/PartRem[18][3] ), .B(
        \u_div/SumTmp[17][3] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_18_3  ( .A(\u_div/PartRem[19][3] ), .B(
        \u_div/SumTmp[18][3] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_19_3  ( .A(\u_div/PartRem[20][3] ), .B(
        \u_div/SumTmp[19][3] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_20_3  ( .A(\u_div/PartRem[21][3] ), .B(
        \u_div/SumTmp[20][3] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_21_3  ( .A(\u_div/PartRem[22][3] ), .B(
        \u_div/SumTmp[21][3] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_22_3  ( .A(\u_div/PartRem[23][3] ), .B(
        \u_div/SumTmp[22][3] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_23_3  ( .A(\u_div/PartRem[24][3] ), .B(
        \u_div/SumTmp[23][3] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_24_3  ( .A(\u_div/PartRem[25][3] ), .B(
        \u_div/SumTmp[24][3] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_25_3  ( .A(\u_div/PartRem[26][3] ), .B(
        \u_div/SumTmp[25][3] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_26_3  ( .A(\u_div/PartRem[27][3] ), .B(
        \u_div/SumTmp[26][3] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_27_3  ( .A(\u_div/PartRem[28][3] ), .B(
        \u_div/SumTmp[27][3] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_28_3  ( .A(\u_div/PartRem[29][3] ), .B(
        \u_div/SumTmp[28][3] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_29_3  ( .A(\u_div/PartRem[30][3] ), .B(
        \u_div/SumTmp[29][3] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_30_3  ( .A(\u_div/PartRem[31][3] ), .B(
        \u_div/SumTmp[30][3] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_31_3  ( .A(\u_div/PartRem[32][3] ), .B(
        \u_div/SumTmp[31][3] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_32_3  ( .A(\u_div/PartRem[33][3] ), .B(
        \u_div/SumTmp[32][3] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_33_3  ( .A(\u_div/PartRem[34][3] ), .B(
        \u_div/SumTmp[33][3] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_34_3  ( .A(\u_div/PartRem[35][3] ), .B(
        \u_div/SumTmp[34][3] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_35_3  ( .A(\u_div/PartRem[36][3] ), .B(
        \u_div/SumTmp[35][3] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_36_3  ( .A(\u_div/PartRem[37][3] ), .B(
        \u_div/SumTmp[36][3] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_37_3  ( .A(\u_div/PartRem[38][3] ), .B(
        \u_div/SumTmp[37][3] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_38_3  ( .A(\u_div/PartRem[39][3] ), .B(
        \u_div/SumTmp[38][3] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_39_3  ( .A(\u_div/PartRem[40][3] ), .B(
        \u_div/SumTmp[39][3] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_40_3  ( .A(\u_div/PartRem[41][3] ), .B(
        \u_div/SumTmp[40][3] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_41_3  ( .A(\u_div/PartRem[42][3] ), .B(
        \u_div/SumTmp[41][3] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_42_3  ( .A(\u_div/PartRem[43][3] ), .B(
        \u_div/SumTmp[42][3] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_43_3  ( .A(\u_div/PartRem[44][3] ), .B(
        \u_div/SumTmp[43][3] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_44_3  ( .A(\u_div/PartRem[45][3] ), .B(
        \u_div/SumTmp[44][3] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_45_3  ( .A(\u_div/PartRem[46][3] ), .B(
        \u_div/SumTmp[45][3] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_46_3  ( .A(\u_div/PartRem[47][3] ), .B(
        \u_div/SumTmp[46][3] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_47_3  ( .A(\u_div/PartRem[48][3] ), .B(
        \u_div/SumTmp[47][3] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_48_3  ( .A(\u_div/PartRem[49][3] ), .B(
        \u_div/SumTmp[48][3] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_49_3  ( .A(\u_div/PartRem[50][3] ), .B(
        \u_div/SumTmp[49][3] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_50_3  ( .A(\u_div/PartRem[51][3] ), .B(
        \u_div/SumTmp[50][3] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_51_3  ( .A(\u_div/PartRem[52][3] ), .B(
        \u_div/SumTmp[51][3] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_52_3  ( .A(\u_div/PartRem[53][3] ), .B(
        \u_div/SumTmp[52][3] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_53_3  ( .A(\u_div/PartRem[54][3] ), .B(
        \u_div/SumTmp[53][3] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_54_3  ( .A(\u_div/PartRem[55][3] ), .B(
        \u_div/SumTmp[54][3] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_55_3  ( .A(\u_div/PartRem[56][3] ), .B(
        \u_div/SumTmp[55][3] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_56_3  ( .A(\u_div/PartRem[57][3] ), .B(
        \u_div/SumTmp[56][3] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_57_3  ( .A(\u_div/PartRem[58][3] ), .B(
        \u_div/SumTmp[57][3] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_58_3  ( .A(\u_div/PartRem[59][3] ), .B(
        \u_div/SumTmp[58][3] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][4] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_3  ( .A(\u_div/PartRem[63][0] ), .B(
        \u_div/SumTmp[59][3] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_14_3  ( .A(\u_div/PartRem[15][3] ), .B(
        \u_div/SumTmp[14][3] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_1_4  ( .A(\u_div/PartRem[2][4] ), .B(
        \u_div/SumTmp[1][4] ), .S0(\u_div/CryTmp[1][6] ), .Y(
        \u_div/PartRem[1][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_15_4  ( .A(\u_div/PartRem[16][4] ), .B(
        \u_div/SumTmp[15][4] ), .S0(\u_div/CryTmp[15][6] ), .Y(
        \u_div/PartRem[15][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_16_4  ( .A(\u_div/PartRem[17][4] ), .B(
        \u_div/SumTmp[16][4] ), .S0(\u_div/CryTmp[16][6] ), .Y(
        \u_div/PartRem[16][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_13_4  ( .A(\u_div/PartRem[14][4] ), .B(
        \u_div/SumTmp[13][4] ), .S0(\u_div/CryTmp[13][6] ), .Y(
        \u_div/PartRem[13][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_14_4  ( .A(\u_div/PartRem[15][4] ), .B(
        \u_div/SumTmp[14][4] ), .S0(\u_div/CryTmp[14][6] ), .Y(
        \u_div/PartRem[14][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_17_4  ( .A(\u_div/PartRem[18][4] ), .B(
        \u_div/SumTmp[17][4] ), .S0(\u_div/CryTmp[17][6] ), .Y(
        \u_div/PartRem[17][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_18_4  ( .A(\u_div/PartRem[19][4] ), .B(
        \u_div/SumTmp[18][4] ), .S0(\u_div/CryTmp[18][6] ), .Y(
        \u_div/PartRem[18][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_19_4  ( .A(\u_div/PartRem[20][4] ), .B(
        \u_div/SumTmp[19][4] ), .S0(\u_div/CryTmp[19][6] ), .Y(
        \u_div/PartRem[19][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_20_4  ( .A(\u_div/PartRem[21][4] ), .B(
        \u_div/SumTmp[20][4] ), .S0(\u_div/CryTmp[20][6] ), .Y(
        \u_div/PartRem[20][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_21_4  ( .A(\u_div/PartRem[22][4] ), .B(
        \u_div/SumTmp[21][4] ), .S0(\u_div/CryTmp[21][6] ), .Y(
        \u_div/PartRem[21][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_22_4  ( .A(\u_div/PartRem[23][4] ), .B(
        \u_div/SumTmp[22][4] ), .S0(\u_div/CryTmp[22][6] ), .Y(
        \u_div/PartRem[22][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_23_4  ( .A(\u_div/PartRem[24][4] ), .B(
        \u_div/SumTmp[23][4] ), .S0(\u_div/CryTmp[23][6] ), .Y(
        \u_div/PartRem[23][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_24_4  ( .A(\u_div/PartRem[25][4] ), .B(
        \u_div/SumTmp[24][4] ), .S0(\u_div/CryTmp[24][6] ), .Y(
        \u_div/PartRem[24][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_25_4  ( .A(\u_div/PartRem[26][4] ), .B(
        \u_div/SumTmp[25][4] ), .S0(\u_div/CryTmp[25][6] ), .Y(
        \u_div/PartRem[25][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_26_4  ( .A(\u_div/PartRem[27][4] ), .B(
        \u_div/SumTmp[26][4] ), .S0(\u_div/CryTmp[26][6] ), .Y(
        \u_div/PartRem[26][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_27_4  ( .A(\u_div/PartRem[28][4] ), .B(
        \u_div/SumTmp[27][4] ), .S0(\u_div/CryTmp[27][6] ), .Y(
        \u_div/PartRem[27][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_28_4  ( .A(\u_div/PartRem[29][4] ), .B(
        \u_div/SumTmp[28][4] ), .S0(\u_div/CryTmp[28][6] ), .Y(
        \u_div/PartRem[28][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_29_4  ( .A(\u_div/PartRem[30][4] ), .B(
        \u_div/SumTmp[29][4] ), .S0(\u_div/CryTmp[29][6] ), .Y(
        \u_div/PartRem[29][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_30_4  ( .A(\u_div/PartRem[31][4] ), .B(
        \u_div/SumTmp[30][4] ), .S0(\u_div/CryTmp[30][6] ), .Y(
        \u_div/PartRem[30][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_31_4  ( .A(\u_div/PartRem[32][4] ), .B(
        \u_div/SumTmp[31][4] ), .S0(\u_div/CryTmp[31][6] ), .Y(
        \u_div/PartRem[31][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_32_4  ( .A(\u_div/PartRem[33][4] ), .B(
        \u_div/SumTmp[32][4] ), .S0(\u_div/CryTmp[32][6] ), .Y(
        \u_div/PartRem[32][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_33_4  ( .A(\u_div/PartRem[34][4] ), .B(
        \u_div/SumTmp[33][4] ), .S0(\u_div/CryTmp[33][6] ), .Y(
        \u_div/PartRem[33][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_34_4  ( .A(\u_div/PartRem[35][4] ), .B(
        \u_div/SumTmp[34][4] ), .S0(\u_div/CryTmp[34][6] ), .Y(
        \u_div/PartRem[34][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_35_4  ( .A(\u_div/PartRem[36][4] ), .B(
        \u_div/SumTmp[35][4] ), .S0(\u_div/CryTmp[35][6] ), .Y(
        \u_div/PartRem[35][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_36_4  ( .A(\u_div/PartRem[37][4] ), .B(
        \u_div/SumTmp[36][4] ), .S0(\u_div/CryTmp[36][6] ), .Y(
        \u_div/PartRem[36][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_37_4  ( .A(\u_div/PartRem[38][4] ), .B(
        \u_div/SumTmp[37][4] ), .S0(\u_div/CryTmp[37][6] ), .Y(
        \u_div/PartRem[37][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_38_4  ( .A(\u_div/PartRem[39][4] ), .B(
        \u_div/SumTmp[38][4] ), .S0(\u_div/CryTmp[38][6] ), .Y(
        \u_div/PartRem[38][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_39_4  ( .A(\u_div/PartRem[40][4] ), .B(
        \u_div/SumTmp[39][4] ), .S0(\u_div/CryTmp[39][6] ), .Y(
        \u_div/PartRem[39][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_40_4  ( .A(\u_div/PartRem[41][4] ), .B(
        \u_div/SumTmp[40][4] ), .S0(\u_div/CryTmp[40][6] ), .Y(
        \u_div/PartRem[40][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_41_4  ( .A(\u_div/PartRem[42][4] ), .B(
        \u_div/SumTmp[41][4] ), .S0(\u_div/CryTmp[41][6] ), .Y(
        \u_div/PartRem[41][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_42_4  ( .A(\u_div/PartRem[43][4] ), .B(
        \u_div/SumTmp[42][4] ), .S0(\u_div/CryTmp[42][6] ), .Y(
        \u_div/PartRem[42][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_43_4  ( .A(\u_div/PartRem[44][4] ), .B(
        \u_div/SumTmp[43][4] ), .S0(\u_div/CryTmp[43][6] ), .Y(
        \u_div/PartRem[43][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_44_4  ( .A(\u_div/PartRem[45][4] ), .B(
        \u_div/SumTmp[44][4] ), .S0(\u_div/CryTmp[44][6] ), .Y(
        \u_div/PartRem[44][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_45_4  ( .A(\u_div/PartRem[46][4] ), .B(
        \u_div/SumTmp[45][4] ), .S0(\u_div/CryTmp[45][6] ), .Y(
        \u_div/PartRem[45][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_46_4  ( .A(\u_div/PartRem[47][4] ), .B(
        \u_div/SumTmp[46][4] ), .S0(\u_div/CryTmp[46][6] ), .Y(
        \u_div/PartRem[46][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_47_4  ( .A(\u_div/PartRem[48][4] ), .B(
        \u_div/SumTmp[47][4] ), .S0(\u_div/CryTmp[47][6] ), .Y(
        \u_div/PartRem[47][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_48_4  ( .A(\u_div/PartRem[49][4] ), .B(
        \u_div/SumTmp[48][4] ), .S0(\u_div/CryTmp[48][6] ), .Y(
        \u_div/PartRem[48][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_49_4  ( .A(\u_div/PartRem[50][4] ), .B(
        \u_div/SumTmp[49][4] ), .S0(\u_div/CryTmp[49][6] ), .Y(
        \u_div/PartRem[49][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_50_4  ( .A(\u_div/PartRem[51][4] ), .B(
        \u_div/SumTmp[50][4] ), .S0(\u_div/CryTmp[50][6] ), .Y(
        \u_div/PartRem[50][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_51_4  ( .A(\u_div/PartRem[52][4] ), .B(
        \u_div/SumTmp[51][4] ), .S0(\u_div/CryTmp[51][6] ), .Y(
        \u_div/PartRem[51][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_52_4  ( .A(\u_div/PartRem[53][4] ), .B(
        \u_div/SumTmp[52][4] ), .S0(\u_div/CryTmp[52][6] ), .Y(
        \u_div/PartRem[52][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_53_4  ( .A(\u_div/PartRem[54][4] ), .B(
        \u_div/SumTmp[53][4] ), .S0(\u_div/CryTmp[53][6] ), .Y(
        \u_div/PartRem[53][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_54_4  ( .A(\u_div/PartRem[55][4] ), .B(
        \u_div/SumTmp[54][4] ), .S0(\u_div/CryTmp[54][6] ), .Y(
        \u_div/PartRem[54][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_55_4  ( .A(\u_div/PartRem[56][4] ), .B(
        \u_div/SumTmp[55][4] ), .S0(\u_div/CryTmp[55][6] ), .Y(
        \u_div/PartRem[55][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_56_4  ( .A(\u_div/PartRem[57][4] ), .B(
        \u_div/SumTmp[56][4] ), .S0(\u_div/CryTmp[56][6] ), .Y(
        \u_div/PartRem[56][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_57_4  ( .A(\u_div/PartRem[58][4] ), .B(
        \u_div/SumTmp[57][4] ), .S0(\u_div/CryTmp[57][6] ), .Y(
        \u_div/PartRem[57][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_58_4  ( .A(\u_div/PartRem[59][4] ), .B(
        \u_div/SumTmp[58][4] ), .S0(\u_div/CryTmp[58][6] ), .Y(
        \u_div/PartRem[58][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_59_4  ( .A(\u_div/PartRem[64][0] ), .B(
        \u_div/SumTmp[59][4] ), .S0(\u_div/CryTmp[59][6] ), .Y(
        \u_div/PartRem[59][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_12_4  ( .A(\u_div/PartRem[13][4] ), .B(
        \u_div/SumTmp[12][4] ), .S0(\u_div/CryTmp[12][6] ), .Y(
        \u_div/PartRem[12][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_10_4  ( .A(\u_div/PartRem[11][4] ), .B(
        \u_div/SumTmp[10][4] ), .S0(\u_div/CryTmp[10][6] ), .Y(
        \u_div/PartRem[10][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_11_4  ( .A(\u_div/PartRem[12][4] ), .B(
        \u_div/SumTmp[11][4] ), .S0(\u_div/CryTmp[11][6] ), .Y(
        \u_div/PartRem[11][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_9_4  ( .A(\u_div/PartRem[10][4] ), .B(
        \u_div/SumTmp[9][4] ), .S0(\u_div/CryTmp[9][6] ), .Y(
        \u_div/PartRem[9][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_7_4  ( .A(\u_div/PartRem[8][4] ), .B(
        \u_div/SumTmp[7][4] ), .S0(\u_div/CryTmp[7][6] ), .Y(
        \u_div/PartRem[7][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_8_4  ( .A(\u_div/PartRem[9][4] ), .B(
        \u_div/SumTmp[8][4] ), .S0(\u_div/CryTmp[8][6] ), .Y(
        \u_div/PartRem[8][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_6_4  ( .A(\u_div/PartRem[7][4] ), .B(
        \u_div/SumTmp[6][4] ), .S0(\u_div/CryTmp[6][6] ), .Y(
        \u_div/PartRem[6][5] ) );
  MX2XL \u_div/u_mx_PartRem_1_4_4  ( .A(\u_div/PartRem[5][4] ), .B(
        \u_div/SumTmp[4][4] ), .S0(\u_div/CryTmp[4][6] ), .Y(
        \u_div/PartRem[4][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_5_4  ( .A(\u_div/PartRem[6][4] ), .B(
        \u_div/SumTmp[5][4] ), .S0(\u_div/CryTmp[5][6] ), .Y(
        \u_div/PartRem[5][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_3_4  ( .A(\u_div/PartRem[4][4] ), .B(
        \u_div/SumTmp[3][4] ), .S0(\u_div/CryTmp[3][6] ), .Y(
        \u_div/PartRem[3][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_1_2_4  ( .A(\u_div/PartRem[3][4] ), .B(
        \u_div/SumTmp[2][4] ), .S0(\u_div/CryTmp[2][6] ), .Y(
        \u_div/PartRem[2][5] ) );
  NOR2BX2 U1 ( .AN(\u_div/PartRem[64][0] ), .B(n6), .Y(\u_div/CryTmp[59][6] )
         );
  XOR2XL U2 ( .A(\u_div/CryTmp[59][6] ), .B(n2), .Y(\u_div/QInv[59] ) );
  INVX3 U3 ( .A(n1), .Y(n2) );
  CLKINVX1 U4 ( .A(n4), .Y(n1) );
  MXI2X1 U5 ( .A(\u_div/SumTmp[1][3] ), .B(\u_div/CryTmp[2][6] ), .S0(
        \u_div/CryTmp[1][6] ), .Y(\u_div/PartRem[1][4] ) );
  CLKINVX1 U6 ( .A(\u_div/CryTmp[2][6] ), .Y(\u_div/SumTmp[1][3] ) );
  MXI2X1 U7 ( .A(\u_div/SumTmp[3][3] ), .B(\u_div/CryTmp[4][6] ), .S0(
        \u_div/CryTmp[3][6] ), .Y(\u_div/PartRem[3][4] ) );
  CLKINVX1 U8 ( .A(\u_div/CryTmp[4][6] ), .Y(\u_div/SumTmp[3][3] ) );
  MXI2X1 U9 ( .A(\u_div/SumTmp[2][3] ), .B(\u_div/CryTmp[3][6] ), .S0(
        \u_div/CryTmp[2][6] ), .Y(\u_div/PartRem[2][4] ) );
  CLKINVX1 U10 ( .A(\u_div/CryTmp[3][6] ), .Y(\u_div/SumTmp[2][3] ) );
  MXI2X1 U11 ( .A(\u_div/SumTmp[4][3] ), .B(\u_div/CryTmp[5][6] ), .S0(
        \u_div/CryTmp[4][6] ), .Y(\u_div/PartRem[4][4] ) );
  CLKINVX1 U12 ( .A(\u_div/CryTmp[5][6] ), .Y(\u_div/SumTmp[4][3] ) );
  MXI2X1 U13 ( .A(\u_div/SumTmp[6][3] ), .B(\u_div/CryTmp[7][6] ), .S0(
        \u_div/CryTmp[6][6] ), .Y(\u_div/PartRem[6][4] ) );
  CLKINVX1 U14 ( .A(\u_div/CryTmp[7][6] ), .Y(\u_div/SumTmp[6][3] ) );
  MXI2X1 U15 ( .A(\u_div/SumTmp[5][3] ), .B(\u_div/CryTmp[6][6] ), .S0(
        \u_div/CryTmp[5][6] ), .Y(\u_div/PartRem[5][4] ) );
  CLKINVX1 U16 ( .A(\u_div/CryTmp[6][6] ), .Y(\u_div/SumTmp[5][3] ) );
  MXI2X1 U17 ( .A(\u_div/SumTmp[7][3] ), .B(\u_div/CryTmp[8][6] ), .S0(
        \u_div/CryTmp[7][6] ), .Y(\u_div/PartRem[7][4] ) );
  CLKINVX1 U18 ( .A(\u_div/CryTmp[8][6] ), .Y(\u_div/SumTmp[7][3] ) );
  MXI2X1 U19 ( .A(\u_div/SumTmp[9][3] ), .B(\u_div/CryTmp[10][6] ), .S0(
        \u_div/CryTmp[9][6] ), .Y(\u_div/PartRem[9][4] ) );
  CLKINVX1 U20 ( .A(\u_div/CryTmp[10][6] ), .Y(\u_div/SumTmp[9][3] ) );
  MXI2X1 U21 ( .A(\u_div/SumTmp[8][3] ), .B(\u_div/CryTmp[9][6] ), .S0(
        \u_div/CryTmp[8][6] ), .Y(\u_div/PartRem[8][4] ) );
  CLKINVX1 U22 ( .A(\u_div/CryTmp[9][6] ), .Y(\u_div/SumTmp[8][3] ) );
  MXI2X1 U23 ( .A(\u_div/SumTmp[10][3] ), .B(\u_div/CryTmp[11][6] ), .S0(
        \u_div/CryTmp[10][6] ), .Y(\u_div/PartRem[10][4] ) );
  CLKINVX1 U24 ( .A(\u_div/CryTmp[11][6] ), .Y(\u_div/SumTmp[10][3] ) );
  MXI2X1 U25 ( .A(\u_div/SumTmp[12][3] ), .B(\u_div/CryTmp[13][6] ), .S0(
        \u_div/CryTmp[12][6] ), .Y(\u_div/PartRem[12][4] ) );
  CLKINVX1 U26 ( .A(\u_div/CryTmp[13][6] ), .Y(\u_div/SumTmp[12][3] ) );
  MXI2X1 U27 ( .A(\u_div/SumTmp[11][3] ), .B(\u_div/CryTmp[12][6] ), .S0(
        \u_div/CryTmp[11][6] ), .Y(\u_div/PartRem[11][4] ) );
  CLKINVX1 U28 ( .A(\u_div/CryTmp[12][6] ), .Y(\u_div/SumTmp[11][3] ) );
  MXI2X1 U29 ( .A(\u_div/SumTmp[13][3] ), .B(\u_div/PartRem[14][3] ), .S0(
        \u_div/CryTmp[13][6] ), .Y(\u_div/PartRem[13][4] ) );
  CLKINVX1 U30 ( .A(\u_div/PartRem[14][3] ), .Y(\u_div/SumTmp[13][3] ) );
  MXI2X1 U31 ( .A(\u_div/SumTmp[14][2] ), .B(\u_div/PartRem[15][2] ), .S0(
        \u_div/CryTmp[14][6] ), .Y(\u_div/PartRem[14][3] ) );
  CLKINVX1 U32 ( .A(\u_div/PartRem[15][2] ), .Y(\u_div/SumTmp[14][2] ) );
  MXI2X1 U33 ( .A(n5), .B(\u_div/PartRem[62][0] ), .S0(\u_div/CryTmp[59][6] ), 
        .Y(\u_div/PartRem[59][3] ) );
  CLKINVX1 U34 ( .A(\u_div/PartRem[62][0] ), .Y(n5) );
  MXI2X1 U35 ( .A(\u_div/SumTmp[58][2] ), .B(\u_div/PartRem[59][2] ), .S0(
        \u_div/CryTmp[58][6] ), .Y(\u_div/PartRem[58][3] ) );
  CLKINVX1 U36 ( .A(\u_div/PartRem[59][2] ), .Y(\u_div/SumTmp[58][2] ) );
  MXI2X1 U37 ( .A(\u_div/SumTmp[57][2] ), .B(\u_div/PartRem[58][2] ), .S0(
        \u_div/CryTmp[57][6] ), .Y(\u_div/PartRem[57][3] ) );
  CLKINVX1 U38 ( .A(\u_div/PartRem[58][2] ), .Y(\u_div/SumTmp[57][2] ) );
  MXI2X1 U39 ( .A(\u_div/SumTmp[56][2] ), .B(\u_div/PartRem[57][2] ), .S0(
        \u_div/CryTmp[56][6] ), .Y(\u_div/PartRem[56][3] ) );
  CLKINVX1 U40 ( .A(\u_div/PartRem[57][2] ), .Y(\u_div/SumTmp[56][2] ) );
  MXI2X1 U41 ( .A(\u_div/SumTmp[55][2] ), .B(\u_div/PartRem[56][2] ), .S0(
        \u_div/CryTmp[55][6] ), .Y(\u_div/PartRem[55][3] ) );
  CLKINVX1 U42 ( .A(\u_div/PartRem[56][2] ), .Y(\u_div/SumTmp[55][2] ) );
  MXI2X1 U43 ( .A(\u_div/SumTmp[54][2] ), .B(\u_div/PartRem[55][2] ), .S0(
        \u_div/CryTmp[54][6] ), .Y(\u_div/PartRem[54][3] ) );
  CLKINVX1 U44 ( .A(\u_div/PartRem[55][2] ), .Y(\u_div/SumTmp[54][2] ) );
  MXI2X1 U45 ( .A(\u_div/SumTmp[53][2] ), .B(\u_div/PartRem[54][2] ), .S0(
        \u_div/CryTmp[53][6] ), .Y(\u_div/PartRem[53][3] ) );
  CLKINVX1 U46 ( .A(\u_div/PartRem[54][2] ), .Y(\u_div/SumTmp[53][2] ) );
  MXI2X1 U47 ( .A(\u_div/SumTmp[52][2] ), .B(\u_div/PartRem[53][2] ), .S0(
        \u_div/CryTmp[52][6] ), .Y(\u_div/PartRem[52][3] ) );
  CLKINVX1 U48 ( .A(\u_div/PartRem[53][2] ), .Y(\u_div/SumTmp[52][2] ) );
  MXI2X1 U49 ( .A(\u_div/SumTmp[51][2] ), .B(\u_div/PartRem[52][2] ), .S0(
        \u_div/CryTmp[51][6] ), .Y(\u_div/PartRem[51][3] ) );
  CLKINVX1 U50 ( .A(\u_div/PartRem[52][2] ), .Y(\u_div/SumTmp[51][2] ) );
  MXI2X1 U51 ( .A(\u_div/SumTmp[50][2] ), .B(\u_div/PartRem[51][2] ), .S0(
        \u_div/CryTmp[50][6] ), .Y(\u_div/PartRem[50][3] ) );
  CLKINVX1 U52 ( .A(\u_div/PartRem[51][2] ), .Y(\u_div/SumTmp[50][2] ) );
  MXI2X1 U53 ( .A(\u_div/SumTmp[49][2] ), .B(\u_div/PartRem[50][2] ), .S0(
        \u_div/CryTmp[49][6] ), .Y(\u_div/PartRem[49][3] ) );
  CLKINVX1 U54 ( .A(\u_div/PartRem[50][2] ), .Y(\u_div/SumTmp[49][2] ) );
  MXI2X1 U55 ( .A(\u_div/SumTmp[48][2] ), .B(\u_div/PartRem[49][2] ), .S0(
        \u_div/CryTmp[48][6] ), .Y(\u_div/PartRem[48][3] ) );
  CLKINVX1 U56 ( .A(\u_div/PartRem[49][2] ), .Y(\u_div/SumTmp[48][2] ) );
  MXI2X1 U57 ( .A(\u_div/SumTmp[47][2] ), .B(\u_div/PartRem[48][2] ), .S0(
        \u_div/CryTmp[47][6] ), .Y(\u_div/PartRem[47][3] ) );
  CLKINVX1 U58 ( .A(\u_div/PartRem[48][2] ), .Y(\u_div/SumTmp[47][2] ) );
  MXI2X1 U59 ( .A(\u_div/SumTmp[46][2] ), .B(\u_div/PartRem[47][2] ), .S0(
        \u_div/CryTmp[46][6] ), .Y(\u_div/PartRem[46][3] ) );
  CLKINVX1 U60 ( .A(\u_div/PartRem[47][2] ), .Y(\u_div/SumTmp[46][2] ) );
  MXI2X1 U61 ( .A(\u_div/SumTmp[45][2] ), .B(\u_div/PartRem[46][2] ), .S0(
        \u_div/CryTmp[45][6] ), .Y(\u_div/PartRem[45][3] ) );
  CLKINVX1 U62 ( .A(\u_div/PartRem[46][2] ), .Y(\u_div/SumTmp[45][2] ) );
  MXI2X1 U63 ( .A(\u_div/SumTmp[44][2] ), .B(\u_div/PartRem[45][2] ), .S0(
        \u_div/CryTmp[44][6] ), .Y(\u_div/PartRem[44][3] ) );
  CLKINVX1 U64 ( .A(\u_div/PartRem[45][2] ), .Y(\u_div/SumTmp[44][2] ) );
  MXI2X1 U65 ( .A(\u_div/SumTmp[43][2] ), .B(\u_div/PartRem[44][2] ), .S0(
        \u_div/CryTmp[43][6] ), .Y(\u_div/PartRem[43][3] ) );
  CLKINVX1 U66 ( .A(\u_div/PartRem[44][2] ), .Y(\u_div/SumTmp[43][2] ) );
  MXI2X1 U67 ( .A(\u_div/SumTmp[42][2] ), .B(\u_div/PartRem[43][2] ), .S0(
        \u_div/CryTmp[42][6] ), .Y(\u_div/PartRem[42][3] ) );
  CLKINVX1 U68 ( .A(\u_div/PartRem[43][2] ), .Y(\u_div/SumTmp[42][2] ) );
  MXI2X1 U69 ( .A(\u_div/SumTmp[41][2] ), .B(\u_div/PartRem[42][2] ), .S0(
        \u_div/CryTmp[41][6] ), .Y(\u_div/PartRem[41][3] ) );
  CLKINVX1 U70 ( .A(\u_div/PartRem[42][2] ), .Y(\u_div/SumTmp[41][2] ) );
  MXI2X1 U71 ( .A(\u_div/SumTmp[40][2] ), .B(\u_div/PartRem[41][2] ), .S0(
        \u_div/CryTmp[40][6] ), .Y(\u_div/PartRem[40][3] ) );
  CLKINVX1 U72 ( .A(\u_div/PartRem[41][2] ), .Y(\u_div/SumTmp[40][2] ) );
  MXI2X1 U73 ( .A(\u_div/SumTmp[39][2] ), .B(\u_div/PartRem[40][2] ), .S0(
        \u_div/CryTmp[39][6] ), .Y(\u_div/PartRem[39][3] ) );
  CLKINVX1 U74 ( .A(\u_div/PartRem[40][2] ), .Y(\u_div/SumTmp[39][2] ) );
  MXI2X1 U75 ( .A(\u_div/SumTmp[38][2] ), .B(\u_div/PartRem[39][2] ), .S0(
        \u_div/CryTmp[38][6] ), .Y(\u_div/PartRem[38][3] ) );
  CLKINVX1 U76 ( .A(\u_div/PartRem[39][2] ), .Y(\u_div/SumTmp[38][2] ) );
  MXI2X1 U77 ( .A(\u_div/SumTmp[37][2] ), .B(\u_div/PartRem[38][2] ), .S0(
        \u_div/CryTmp[37][6] ), .Y(\u_div/PartRem[37][3] ) );
  CLKINVX1 U78 ( .A(\u_div/PartRem[38][2] ), .Y(\u_div/SumTmp[37][2] ) );
  MXI2X1 U79 ( .A(\u_div/SumTmp[36][2] ), .B(\u_div/PartRem[37][2] ), .S0(
        \u_div/CryTmp[36][6] ), .Y(\u_div/PartRem[36][3] ) );
  CLKINVX1 U80 ( .A(\u_div/PartRem[37][2] ), .Y(\u_div/SumTmp[36][2] ) );
  MXI2X1 U81 ( .A(\u_div/SumTmp[35][2] ), .B(\u_div/PartRem[36][2] ), .S0(
        \u_div/CryTmp[35][6] ), .Y(\u_div/PartRem[35][3] ) );
  CLKINVX1 U82 ( .A(\u_div/PartRem[36][2] ), .Y(\u_div/SumTmp[35][2] ) );
  MXI2X1 U83 ( .A(\u_div/SumTmp[34][2] ), .B(\u_div/PartRem[35][2] ), .S0(
        \u_div/CryTmp[34][6] ), .Y(\u_div/PartRem[34][3] ) );
  CLKINVX1 U84 ( .A(\u_div/PartRem[35][2] ), .Y(\u_div/SumTmp[34][2] ) );
  MXI2X1 U85 ( .A(\u_div/SumTmp[33][2] ), .B(\u_div/PartRem[34][2] ), .S0(
        \u_div/CryTmp[33][6] ), .Y(\u_div/PartRem[33][3] ) );
  CLKINVX1 U86 ( .A(\u_div/PartRem[34][2] ), .Y(\u_div/SumTmp[33][2] ) );
  MXI2X1 U87 ( .A(\u_div/SumTmp[32][2] ), .B(\u_div/PartRem[33][2] ), .S0(
        \u_div/CryTmp[32][6] ), .Y(\u_div/PartRem[32][3] ) );
  CLKINVX1 U88 ( .A(\u_div/PartRem[33][2] ), .Y(\u_div/SumTmp[32][2] ) );
  MXI2X1 U89 ( .A(\u_div/SumTmp[31][2] ), .B(\u_div/PartRem[32][2] ), .S0(
        \u_div/CryTmp[31][6] ), .Y(\u_div/PartRem[31][3] ) );
  CLKINVX1 U90 ( .A(\u_div/PartRem[32][2] ), .Y(\u_div/SumTmp[31][2] ) );
  MXI2X1 U91 ( .A(\u_div/SumTmp[30][2] ), .B(\u_div/PartRem[31][2] ), .S0(
        \u_div/CryTmp[30][6] ), .Y(\u_div/PartRem[30][3] ) );
  CLKINVX1 U92 ( .A(\u_div/PartRem[31][2] ), .Y(\u_div/SumTmp[30][2] ) );
  MXI2X1 U93 ( .A(\u_div/SumTmp[29][2] ), .B(\u_div/PartRem[30][2] ), .S0(
        \u_div/CryTmp[29][6] ), .Y(\u_div/PartRem[29][3] ) );
  CLKINVX1 U94 ( .A(\u_div/PartRem[30][2] ), .Y(\u_div/SumTmp[29][2] ) );
  MXI2X1 U95 ( .A(\u_div/SumTmp[28][2] ), .B(\u_div/PartRem[29][2] ), .S0(
        \u_div/CryTmp[28][6] ), .Y(\u_div/PartRem[28][3] ) );
  CLKINVX1 U96 ( .A(\u_div/PartRem[29][2] ), .Y(\u_div/SumTmp[28][2] ) );
  MXI2X1 U97 ( .A(\u_div/SumTmp[27][2] ), .B(\u_div/PartRem[28][2] ), .S0(
        \u_div/CryTmp[27][6] ), .Y(\u_div/PartRem[27][3] ) );
  CLKINVX1 U98 ( .A(\u_div/PartRem[28][2] ), .Y(\u_div/SumTmp[27][2] ) );
  MXI2X1 U99 ( .A(\u_div/SumTmp[26][2] ), .B(\u_div/PartRem[27][2] ), .S0(
        \u_div/CryTmp[26][6] ), .Y(\u_div/PartRem[26][3] ) );
  CLKINVX1 U100 ( .A(\u_div/PartRem[27][2] ), .Y(\u_div/SumTmp[26][2] ) );
  MXI2X1 U101 ( .A(\u_div/SumTmp[25][2] ), .B(\u_div/PartRem[26][2] ), .S0(
        \u_div/CryTmp[25][6] ), .Y(\u_div/PartRem[25][3] ) );
  CLKINVX1 U102 ( .A(\u_div/PartRem[26][2] ), .Y(\u_div/SumTmp[25][2] ) );
  MXI2X1 U103 ( .A(\u_div/SumTmp[24][2] ), .B(\u_div/PartRem[25][2] ), .S0(
        \u_div/CryTmp[24][6] ), .Y(\u_div/PartRem[24][3] ) );
  CLKINVX1 U104 ( .A(\u_div/PartRem[25][2] ), .Y(\u_div/SumTmp[24][2] ) );
  MXI2X1 U105 ( .A(\u_div/SumTmp[23][2] ), .B(\u_div/PartRem[24][2] ), .S0(
        \u_div/CryTmp[23][6] ), .Y(\u_div/PartRem[23][3] ) );
  CLKINVX1 U106 ( .A(\u_div/PartRem[24][2] ), .Y(\u_div/SumTmp[23][2] ) );
  MXI2X1 U107 ( .A(\u_div/SumTmp[22][2] ), .B(\u_div/PartRem[23][2] ), .S0(
        \u_div/CryTmp[22][6] ), .Y(\u_div/PartRem[22][3] ) );
  CLKINVX1 U108 ( .A(\u_div/PartRem[23][2] ), .Y(\u_div/SumTmp[22][2] ) );
  MXI2X1 U109 ( .A(\u_div/SumTmp[21][2] ), .B(\u_div/PartRem[22][2] ), .S0(
        \u_div/CryTmp[21][6] ), .Y(\u_div/PartRem[21][3] ) );
  CLKINVX1 U110 ( .A(\u_div/PartRem[22][2] ), .Y(\u_div/SumTmp[21][2] ) );
  MXI2X1 U111 ( .A(\u_div/SumTmp[20][2] ), .B(\u_div/PartRem[21][2] ), .S0(
        \u_div/CryTmp[20][6] ), .Y(\u_div/PartRem[20][3] ) );
  CLKINVX1 U112 ( .A(\u_div/PartRem[21][2] ), .Y(\u_div/SumTmp[20][2] ) );
  MXI2X1 U113 ( .A(\u_div/SumTmp[19][2] ), .B(\u_div/PartRem[20][2] ), .S0(
        \u_div/CryTmp[19][6] ), .Y(\u_div/PartRem[19][3] ) );
  CLKINVX1 U114 ( .A(\u_div/PartRem[20][2] ), .Y(\u_div/SumTmp[19][2] ) );
  MXI2X1 U115 ( .A(\u_div/SumTmp[18][2] ), .B(\u_div/PartRem[19][2] ), .S0(
        \u_div/CryTmp[18][6] ), .Y(\u_div/PartRem[18][3] ) );
  CLKINVX1 U116 ( .A(\u_div/PartRem[19][2] ), .Y(\u_div/SumTmp[18][2] ) );
  MXI2X1 U117 ( .A(\u_div/SumTmp[17][2] ), .B(\u_div/PartRem[18][2] ), .S0(
        \u_div/CryTmp[17][6] ), .Y(\u_div/PartRem[17][3] ) );
  CLKINVX1 U118 ( .A(\u_div/PartRem[18][2] ), .Y(\u_div/SumTmp[17][2] ) );
  MXI2X1 U119 ( .A(\u_div/SumTmp[16][2] ), .B(\u_div/PartRem[17][2] ), .S0(
        \u_div/CryTmp[16][6] ), .Y(\u_div/PartRem[16][3] ) );
  CLKINVX1 U120 ( .A(\u_div/PartRem[17][2] ), .Y(\u_div/SumTmp[16][2] ) );
  MXI2X1 U121 ( .A(\u_div/SumTmp[15][2] ), .B(\u_div/PartRem[16][2] ), .S0(
        \u_div/CryTmp[15][6] ), .Y(\u_div/PartRem[15][3] ) );
  CLKINVX1 U122 ( .A(\u_div/PartRem[16][2] ), .Y(\u_div/SumTmp[15][2] ) );
  INVX4 U123 ( .A(n1), .Y(n3) );
  CLKBUFX3 U124 ( .A(\u_div/QInv[63] ), .Y(n4) );
  OR2X1 U125 ( .A(\u_div/PartRem[59][5] ), .B(\u_div/u_add_PartRem_2_58/n2 ), 
        .Y(\u_div/CryTmp[58][6] ) );
  XNOR2X1 U126 ( .A(\u_div/PartRem[59][3] ), .B(\u_div/PartRem[59][2] ), .Y(
        \u_div/SumTmp[58][3] ) );
  OR2X1 U127 ( .A(\u_div/PartRem[59][2] ), .B(\u_div/PartRem[59][3] ), .Y(
        \u_div/u_add_PartRem_2_58/n3 ) );
  OR2X1 U128 ( .A(\u_div/PartRem[58][5] ), .B(\u_div/u_add_PartRem_2_57/n2 ), 
        .Y(\u_div/CryTmp[57][6] ) );
  XNOR2X1 U129 ( .A(\u_div/PartRem[58][3] ), .B(\u_div/PartRem[58][2] ), .Y(
        \u_div/SumTmp[57][3] ) );
  OR2X1 U130 ( .A(\u_div/PartRem[58][2] ), .B(\u_div/PartRem[58][3] ), .Y(
        \u_div/u_add_PartRem_2_57/n3 ) );
  OR2X1 U131 ( .A(\u_div/PartRem[57][5] ), .B(\u_div/u_add_PartRem_2_56/n2 ), 
        .Y(\u_div/CryTmp[56][6] ) );
  XNOR2X1 U132 ( .A(\u_div/PartRem[57][3] ), .B(\u_div/PartRem[57][2] ), .Y(
        \u_div/SumTmp[56][3] ) );
  OR2X1 U133 ( .A(\u_div/PartRem[57][2] ), .B(\u_div/PartRem[57][3] ), .Y(
        \u_div/u_add_PartRem_2_56/n3 ) );
  OR2X1 U134 ( .A(\u_div/PartRem[56][5] ), .B(\u_div/u_add_PartRem_2_55/n2 ), 
        .Y(\u_div/CryTmp[55][6] ) );
  XNOR2X1 U135 ( .A(\u_div/PartRem[56][3] ), .B(\u_div/PartRem[56][2] ), .Y(
        \u_div/SumTmp[55][3] ) );
  OR2X1 U136 ( .A(\u_div/PartRem[56][2] ), .B(\u_div/PartRem[56][3] ), .Y(
        \u_div/u_add_PartRem_2_55/n3 ) );
  OR2X1 U137 ( .A(\u_div/PartRem[55][5] ), .B(\u_div/u_add_PartRem_2_54/n2 ), 
        .Y(\u_div/CryTmp[54][6] ) );
  XNOR2X1 U138 ( .A(\u_div/PartRem[55][3] ), .B(\u_div/PartRem[55][2] ), .Y(
        \u_div/SumTmp[54][3] ) );
  OR2X1 U139 ( .A(\u_div/PartRem[55][2] ), .B(\u_div/PartRem[55][3] ), .Y(
        \u_div/u_add_PartRem_2_54/n3 ) );
  OR2X1 U140 ( .A(\u_div/PartRem[54][5] ), .B(\u_div/u_add_PartRem_2_53/n2 ), 
        .Y(\u_div/CryTmp[53][6] ) );
  XNOR2X1 U141 ( .A(\u_div/PartRem[54][3] ), .B(\u_div/PartRem[54][2] ), .Y(
        \u_div/SumTmp[53][3] ) );
  OR2X1 U142 ( .A(\u_div/PartRem[54][2] ), .B(\u_div/PartRem[54][3] ), .Y(
        \u_div/u_add_PartRem_2_53/n3 ) );
  OR2X1 U143 ( .A(\u_div/PartRem[53][5] ), .B(\u_div/u_add_PartRem_2_52/n2 ), 
        .Y(\u_div/CryTmp[52][6] ) );
  XNOR2X1 U144 ( .A(\u_div/PartRem[53][3] ), .B(\u_div/PartRem[53][2] ), .Y(
        \u_div/SumTmp[52][3] ) );
  OR2X1 U145 ( .A(\u_div/PartRem[53][2] ), .B(\u_div/PartRem[53][3] ), .Y(
        \u_div/u_add_PartRem_2_52/n3 ) );
  OR2X1 U146 ( .A(\u_div/PartRem[52][5] ), .B(\u_div/u_add_PartRem_2_51/n2 ), 
        .Y(\u_div/CryTmp[51][6] ) );
  XNOR2X1 U147 ( .A(\u_div/PartRem[52][3] ), .B(\u_div/PartRem[52][2] ), .Y(
        \u_div/SumTmp[51][3] ) );
  OR2X1 U148 ( .A(\u_div/PartRem[52][2] ), .B(\u_div/PartRem[52][3] ), .Y(
        \u_div/u_add_PartRem_2_51/n3 ) );
  OR2X1 U149 ( .A(\u_div/PartRem[51][5] ), .B(\u_div/u_add_PartRem_2_50/n2 ), 
        .Y(\u_div/CryTmp[50][6] ) );
  XNOR2X1 U150 ( .A(\u_div/PartRem[51][3] ), .B(\u_div/PartRem[51][2] ), .Y(
        \u_div/SumTmp[50][3] ) );
  OR2X1 U151 ( .A(\u_div/PartRem[51][2] ), .B(\u_div/PartRem[51][3] ), .Y(
        \u_div/u_add_PartRem_2_50/n3 ) );
  OR2X1 U152 ( .A(\u_div/PartRem[50][5] ), .B(\u_div/u_add_PartRem_2_49/n2 ), 
        .Y(\u_div/CryTmp[49][6] ) );
  XNOR2X1 U153 ( .A(\u_div/PartRem[50][3] ), .B(\u_div/PartRem[50][2] ), .Y(
        \u_div/SumTmp[49][3] ) );
  OR2X1 U154 ( .A(\u_div/PartRem[50][2] ), .B(\u_div/PartRem[50][3] ), .Y(
        \u_div/u_add_PartRem_2_49/n3 ) );
  OR2X1 U155 ( .A(\u_div/PartRem[49][5] ), .B(\u_div/u_add_PartRem_2_48/n2 ), 
        .Y(\u_div/CryTmp[48][6] ) );
  XNOR2X1 U156 ( .A(\u_div/PartRem[49][3] ), .B(\u_div/PartRem[49][2] ), .Y(
        \u_div/SumTmp[48][3] ) );
  OR2X1 U157 ( .A(\u_div/PartRem[49][2] ), .B(\u_div/PartRem[49][3] ), .Y(
        \u_div/u_add_PartRem_2_48/n3 ) );
  OR2X1 U158 ( .A(\u_div/PartRem[48][5] ), .B(\u_div/u_add_PartRem_2_47/n2 ), 
        .Y(\u_div/CryTmp[47][6] ) );
  XNOR2X1 U159 ( .A(\u_div/PartRem[48][3] ), .B(\u_div/PartRem[48][2] ), .Y(
        \u_div/SumTmp[47][3] ) );
  OR2X1 U160 ( .A(\u_div/PartRem[48][2] ), .B(\u_div/PartRem[48][3] ), .Y(
        \u_div/u_add_PartRem_2_47/n3 ) );
  OR2X1 U161 ( .A(\u_div/PartRem[47][5] ), .B(\u_div/u_add_PartRem_2_46/n2 ), 
        .Y(\u_div/CryTmp[46][6] ) );
  XNOR2X1 U162 ( .A(\u_div/PartRem[47][3] ), .B(\u_div/PartRem[47][2] ), .Y(
        \u_div/SumTmp[46][3] ) );
  OR2X1 U163 ( .A(\u_div/PartRem[47][2] ), .B(\u_div/PartRem[47][3] ), .Y(
        \u_div/u_add_PartRem_2_46/n3 ) );
  OR2X1 U164 ( .A(\u_div/PartRem[46][5] ), .B(\u_div/u_add_PartRem_2_45/n2 ), 
        .Y(\u_div/CryTmp[45][6] ) );
  XNOR2X1 U165 ( .A(\u_div/PartRem[46][3] ), .B(\u_div/PartRem[46][2] ), .Y(
        \u_div/SumTmp[45][3] ) );
  OR2X1 U166 ( .A(\u_div/PartRem[46][2] ), .B(\u_div/PartRem[46][3] ), .Y(
        \u_div/u_add_PartRem_2_45/n3 ) );
  OR2X1 U167 ( .A(\u_div/PartRem[45][5] ), .B(\u_div/u_add_PartRem_2_44/n2 ), 
        .Y(\u_div/CryTmp[44][6] ) );
  XNOR2X1 U168 ( .A(\u_div/PartRem[45][3] ), .B(\u_div/PartRem[45][2] ), .Y(
        \u_div/SumTmp[44][3] ) );
  OR2X1 U169 ( .A(\u_div/PartRem[45][2] ), .B(\u_div/PartRem[45][3] ), .Y(
        \u_div/u_add_PartRem_2_44/n3 ) );
  OR2X1 U170 ( .A(\u_div/PartRem[44][5] ), .B(\u_div/u_add_PartRem_2_43/n2 ), 
        .Y(\u_div/CryTmp[43][6] ) );
  XNOR2X1 U171 ( .A(\u_div/PartRem[44][3] ), .B(\u_div/PartRem[44][2] ), .Y(
        \u_div/SumTmp[43][3] ) );
  OR2X1 U172 ( .A(\u_div/PartRem[44][2] ), .B(\u_div/PartRem[44][3] ), .Y(
        \u_div/u_add_PartRem_2_43/n3 ) );
  OR2X1 U173 ( .A(\u_div/PartRem[43][5] ), .B(\u_div/u_add_PartRem_2_42/n2 ), 
        .Y(\u_div/CryTmp[42][6] ) );
  XNOR2X1 U174 ( .A(\u_div/PartRem[43][3] ), .B(\u_div/PartRem[43][2] ), .Y(
        \u_div/SumTmp[42][3] ) );
  OR2X1 U175 ( .A(\u_div/PartRem[43][2] ), .B(\u_div/PartRem[43][3] ), .Y(
        \u_div/u_add_PartRem_2_42/n3 ) );
  OR2X1 U176 ( .A(\u_div/PartRem[42][5] ), .B(\u_div/u_add_PartRem_2_41/n2 ), 
        .Y(\u_div/CryTmp[41][6] ) );
  XNOR2X1 U177 ( .A(\u_div/PartRem[42][3] ), .B(\u_div/PartRem[42][2] ), .Y(
        \u_div/SumTmp[41][3] ) );
  OR2X1 U178 ( .A(\u_div/PartRem[42][2] ), .B(\u_div/PartRem[42][3] ), .Y(
        \u_div/u_add_PartRem_2_41/n3 ) );
  OR2X1 U179 ( .A(\u_div/PartRem[41][5] ), .B(\u_div/u_add_PartRem_2_40/n2 ), 
        .Y(\u_div/CryTmp[40][6] ) );
  XNOR2X1 U180 ( .A(\u_div/PartRem[41][3] ), .B(\u_div/PartRem[41][2] ), .Y(
        \u_div/SumTmp[40][3] ) );
  OR2X1 U181 ( .A(\u_div/PartRem[41][2] ), .B(\u_div/PartRem[41][3] ), .Y(
        \u_div/u_add_PartRem_2_40/n3 ) );
  OR2X1 U182 ( .A(\u_div/PartRem[40][5] ), .B(\u_div/u_add_PartRem_2_39/n2 ), 
        .Y(\u_div/CryTmp[39][6] ) );
  XNOR2X1 U183 ( .A(\u_div/PartRem[40][3] ), .B(\u_div/PartRem[40][2] ), .Y(
        \u_div/SumTmp[39][3] ) );
  OR2X1 U184 ( .A(\u_div/PartRem[40][2] ), .B(\u_div/PartRem[40][3] ), .Y(
        \u_div/u_add_PartRem_2_39/n3 ) );
  OR2X1 U185 ( .A(\u_div/PartRem[39][5] ), .B(\u_div/u_add_PartRem_2_38/n2 ), 
        .Y(\u_div/CryTmp[38][6] ) );
  XNOR2X1 U186 ( .A(\u_div/PartRem[39][3] ), .B(\u_div/PartRem[39][2] ), .Y(
        \u_div/SumTmp[38][3] ) );
  OR2X1 U187 ( .A(\u_div/PartRem[39][2] ), .B(\u_div/PartRem[39][3] ), .Y(
        \u_div/u_add_PartRem_2_38/n3 ) );
  OR2X1 U188 ( .A(\u_div/PartRem[38][5] ), .B(\u_div/u_add_PartRem_2_37/n2 ), 
        .Y(\u_div/CryTmp[37][6] ) );
  XNOR2X1 U189 ( .A(\u_div/PartRem[38][3] ), .B(\u_div/PartRem[38][2] ), .Y(
        \u_div/SumTmp[37][3] ) );
  OR2X1 U190 ( .A(\u_div/PartRem[38][2] ), .B(\u_div/PartRem[38][3] ), .Y(
        \u_div/u_add_PartRem_2_37/n3 ) );
  OR2X1 U191 ( .A(\u_div/PartRem[37][5] ), .B(\u_div/u_add_PartRem_2_36/n2 ), 
        .Y(\u_div/CryTmp[36][6] ) );
  XNOR2X1 U192 ( .A(\u_div/PartRem[37][3] ), .B(\u_div/PartRem[37][2] ), .Y(
        \u_div/SumTmp[36][3] ) );
  OR2X1 U193 ( .A(\u_div/PartRem[37][2] ), .B(\u_div/PartRem[37][3] ), .Y(
        \u_div/u_add_PartRem_2_36/n3 ) );
  OR2X1 U194 ( .A(\u_div/PartRem[36][5] ), .B(\u_div/u_add_PartRem_2_35/n2 ), 
        .Y(\u_div/CryTmp[35][6] ) );
  XNOR2X1 U195 ( .A(\u_div/PartRem[36][3] ), .B(\u_div/PartRem[36][2] ), .Y(
        \u_div/SumTmp[35][3] ) );
  OR2X1 U196 ( .A(\u_div/PartRem[36][2] ), .B(\u_div/PartRem[36][3] ), .Y(
        \u_div/u_add_PartRem_2_35/n3 ) );
  OR2X1 U197 ( .A(\u_div/PartRem[35][5] ), .B(\u_div/u_add_PartRem_2_34/n2 ), 
        .Y(\u_div/CryTmp[34][6] ) );
  XNOR2X1 U198 ( .A(\u_div/PartRem[35][3] ), .B(\u_div/PartRem[35][2] ), .Y(
        \u_div/SumTmp[34][3] ) );
  OR2X1 U199 ( .A(\u_div/PartRem[35][2] ), .B(\u_div/PartRem[35][3] ), .Y(
        \u_div/u_add_PartRem_2_34/n3 ) );
  OR2X1 U200 ( .A(\u_div/PartRem[34][5] ), .B(\u_div/u_add_PartRem_2_33/n2 ), 
        .Y(\u_div/CryTmp[33][6] ) );
  XNOR2X1 U201 ( .A(\u_div/PartRem[34][3] ), .B(\u_div/PartRem[34][2] ), .Y(
        \u_div/SumTmp[33][3] ) );
  OR2X1 U202 ( .A(\u_div/PartRem[34][2] ), .B(\u_div/PartRem[34][3] ), .Y(
        \u_div/u_add_PartRem_2_33/n3 ) );
  OR2X1 U203 ( .A(\u_div/PartRem[33][5] ), .B(\u_div/u_add_PartRem_2_32/n2 ), 
        .Y(\u_div/CryTmp[32][6] ) );
  XNOR2X1 U204 ( .A(\u_div/PartRem[33][3] ), .B(\u_div/PartRem[33][2] ), .Y(
        \u_div/SumTmp[32][3] ) );
  OR2X1 U205 ( .A(\u_div/PartRem[33][2] ), .B(\u_div/PartRem[33][3] ), .Y(
        \u_div/u_add_PartRem_2_32/n3 ) );
  OR2X1 U206 ( .A(\u_div/PartRem[32][5] ), .B(\u_div/u_add_PartRem_2_31/n2 ), 
        .Y(\u_div/CryTmp[31][6] ) );
  XNOR2X1 U207 ( .A(\u_div/PartRem[32][3] ), .B(\u_div/PartRem[32][2] ), .Y(
        \u_div/SumTmp[31][3] ) );
  OR2X1 U208 ( .A(\u_div/PartRem[32][2] ), .B(\u_div/PartRem[32][3] ), .Y(
        \u_div/u_add_PartRem_2_31/n3 ) );
  OR2X1 U209 ( .A(\u_div/PartRem[31][5] ), .B(\u_div/u_add_PartRem_2_30/n2 ), 
        .Y(\u_div/CryTmp[30][6] ) );
  XNOR2X1 U210 ( .A(\u_div/PartRem[31][3] ), .B(\u_div/PartRem[31][2] ), .Y(
        \u_div/SumTmp[30][3] ) );
  OR2X1 U211 ( .A(\u_div/PartRem[31][2] ), .B(\u_div/PartRem[31][3] ), .Y(
        \u_div/u_add_PartRem_2_30/n3 ) );
  OR2X1 U212 ( .A(\u_div/PartRem[30][5] ), .B(\u_div/u_add_PartRem_2_29/n2 ), 
        .Y(\u_div/CryTmp[29][6] ) );
  XNOR2X1 U213 ( .A(\u_div/PartRem[30][3] ), .B(\u_div/PartRem[30][2] ), .Y(
        \u_div/SumTmp[29][3] ) );
  OR2X1 U214 ( .A(\u_div/PartRem[30][2] ), .B(\u_div/PartRem[30][3] ), .Y(
        \u_div/u_add_PartRem_2_29/n3 ) );
  OR2X1 U215 ( .A(\u_div/PartRem[29][5] ), .B(\u_div/u_add_PartRem_2_28/n2 ), 
        .Y(\u_div/CryTmp[28][6] ) );
  XNOR2X1 U216 ( .A(\u_div/PartRem[29][3] ), .B(\u_div/PartRem[29][2] ), .Y(
        \u_div/SumTmp[28][3] ) );
  OR2X1 U217 ( .A(\u_div/PartRem[29][2] ), .B(\u_div/PartRem[29][3] ), .Y(
        \u_div/u_add_PartRem_2_28/n3 ) );
  OR2X1 U218 ( .A(\u_div/PartRem[28][5] ), .B(\u_div/u_add_PartRem_2_27/n2 ), 
        .Y(\u_div/CryTmp[27][6] ) );
  XNOR2X1 U219 ( .A(\u_div/PartRem[28][3] ), .B(\u_div/PartRem[28][2] ), .Y(
        \u_div/SumTmp[27][3] ) );
  OR2X1 U220 ( .A(\u_div/PartRem[28][2] ), .B(\u_div/PartRem[28][3] ), .Y(
        \u_div/u_add_PartRem_2_27/n3 ) );
  OR2X1 U221 ( .A(\u_div/PartRem[27][5] ), .B(\u_div/u_add_PartRem_2_26/n2 ), 
        .Y(\u_div/CryTmp[26][6] ) );
  XNOR2X1 U222 ( .A(\u_div/PartRem[27][3] ), .B(\u_div/PartRem[27][2] ), .Y(
        \u_div/SumTmp[26][3] ) );
  OR2X1 U223 ( .A(\u_div/PartRem[27][2] ), .B(\u_div/PartRem[27][3] ), .Y(
        \u_div/u_add_PartRem_2_26/n3 ) );
  OR2X1 U224 ( .A(\u_div/PartRem[26][5] ), .B(\u_div/u_add_PartRem_2_25/n2 ), 
        .Y(\u_div/CryTmp[25][6] ) );
  XNOR2X1 U225 ( .A(\u_div/PartRem[26][3] ), .B(\u_div/PartRem[26][2] ), .Y(
        \u_div/SumTmp[25][3] ) );
  OR2X1 U226 ( .A(\u_div/PartRem[26][2] ), .B(\u_div/PartRem[26][3] ), .Y(
        \u_div/u_add_PartRem_2_25/n3 ) );
  OR2X1 U227 ( .A(\u_div/PartRem[25][5] ), .B(\u_div/u_add_PartRem_2_24/n2 ), 
        .Y(\u_div/CryTmp[24][6] ) );
  XNOR2X1 U228 ( .A(\u_div/PartRem[25][3] ), .B(\u_div/PartRem[25][2] ), .Y(
        \u_div/SumTmp[24][3] ) );
  OR2X1 U229 ( .A(\u_div/PartRem[25][2] ), .B(\u_div/PartRem[25][3] ), .Y(
        \u_div/u_add_PartRem_2_24/n3 ) );
  OR2X1 U230 ( .A(\u_div/PartRem[24][5] ), .B(\u_div/u_add_PartRem_2_23/n2 ), 
        .Y(\u_div/CryTmp[23][6] ) );
  XNOR2X1 U231 ( .A(\u_div/PartRem[24][3] ), .B(\u_div/PartRem[24][2] ), .Y(
        \u_div/SumTmp[23][3] ) );
  OR2X1 U232 ( .A(\u_div/PartRem[24][2] ), .B(\u_div/PartRem[24][3] ), .Y(
        \u_div/u_add_PartRem_2_23/n3 ) );
  OR2X1 U233 ( .A(\u_div/PartRem[23][5] ), .B(\u_div/u_add_PartRem_2_22/n2 ), 
        .Y(\u_div/CryTmp[22][6] ) );
  XNOR2X1 U234 ( .A(\u_div/PartRem[23][3] ), .B(\u_div/PartRem[23][2] ), .Y(
        \u_div/SumTmp[22][3] ) );
  OR2X1 U235 ( .A(\u_div/PartRem[23][2] ), .B(\u_div/PartRem[23][3] ), .Y(
        \u_div/u_add_PartRem_2_22/n3 ) );
  OR2X1 U236 ( .A(\u_div/PartRem[22][5] ), .B(\u_div/u_add_PartRem_2_21/n2 ), 
        .Y(\u_div/CryTmp[21][6] ) );
  XNOR2X1 U237 ( .A(\u_div/PartRem[22][3] ), .B(\u_div/PartRem[22][2] ), .Y(
        \u_div/SumTmp[21][3] ) );
  OR2X1 U238 ( .A(\u_div/PartRem[22][2] ), .B(\u_div/PartRem[22][3] ), .Y(
        \u_div/u_add_PartRem_2_21/n3 ) );
  OR2X1 U239 ( .A(\u_div/PartRem[21][5] ), .B(\u_div/u_add_PartRem_2_20/n2 ), 
        .Y(\u_div/CryTmp[20][6] ) );
  XNOR2X1 U240 ( .A(\u_div/PartRem[21][3] ), .B(\u_div/PartRem[21][2] ), .Y(
        \u_div/SumTmp[20][3] ) );
  OR2X1 U241 ( .A(\u_div/PartRem[21][2] ), .B(\u_div/PartRem[21][3] ), .Y(
        \u_div/u_add_PartRem_2_20/n3 ) );
  OR2X1 U242 ( .A(\u_div/PartRem[20][5] ), .B(\u_div/u_add_PartRem_2_19/n2 ), 
        .Y(\u_div/CryTmp[19][6] ) );
  XNOR2X1 U243 ( .A(\u_div/PartRem[20][3] ), .B(\u_div/PartRem[20][2] ), .Y(
        \u_div/SumTmp[19][3] ) );
  OR2X1 U244 ( .A(\u_div/PartRem[20][2] ), .B(\u_div/PartRem[20][3] ), .Y(
        \u_div/u_add_PartRem_2_19/n3 ) );
  OR2X1 U245 ( .A(\u_div/PartRem[19][5] ), .B(\u_div/u_add_PartRem_2_18/n2 ), 
        .Y(\u_div/CryTmp[18][6] ) );
  XNOR2X1 U246 ( .A(\u_div/PartRem[19][3] ), .B(\u_div/PartRem[19][2] ), .Y(
        \u_div/SumTmp[18][3] ) );
  OR2X1 U247 ( .A(\u_div/PartRem[19][2] ), .B(\u_div/PartRem[19][3] ), .Y(
        \u_div/u_add_PartRem_2_18/n3 ) );
  OR2X1 U248 ( .A(\u_div/PartRem[18][5] ), .B(\u_div/u_add_PartRem_2_17/n2 ), 
        .Y(\u_div/CryTmp[17][6] ) );
  XNOR2X1 U249 ( .A(\u_div/PartRem[18][3] ), .B(\u_div/PartRem[18][2] ), .Y(
        \u_div/SumTmp[17][3] ) );
  OR2X1 U250 ( .A(\u_div/PartRem[18][2] ), .B(\u_div/PartRem[18][3] ), .Y(
        \u_div/u_add_PartRem_2_17/n3 ) );
  OR2X1 U251 ( .A(\u_div/PartRem[17][5] ), .B(\u_div/u_add_PartRem_2_16/n2 ), 
        .Y(\u_div/CryTmp[16][6] ) );
  XNOR2X1 U252 ( .A(\u_div/PartRem[17][3] ), .B(\u_div/PartRem[17][2] ), .Y(
        \u_div/SumTmp[16][3] ) );
  OR2X1 U253 ( .A(\u_div/PartRem[17][2] ), .B(\u_div/PartRem[17][3] ), .Y(
        \u_div/u_add_PartRem_2_16/n3 ) );
  OR2X1 U254 ( .A(\u_div/PartRem[16][5] ), .B(\u_div/u_add_PartRem_2_15/n2 ), 
        .Y(\u_div/CryTmp[15][6] ) );
  XNOR2X1 U255 ( .A(\u_div/PartRem[16][3] ), .B(\u_div/PartRem[16][2] ), .Y(
        \u_div/SumTmp[15][3] ) );
  OR2X1 U256 ( .A(\u_div/PartRem[16][2] ), .B(\u_div/PartRem[16][3] ), .Y(
        \u_div/u_add_PartRem_2_15/n3 ) );
  OR2X1 U257 ( .A(\u_div/PartRem[15][5] ), .B(\u_div/u_add_PartRem_2_14/n2 ), 
        .Y(\u_div/CryTmp[14][6] ) );
  XNOR2X1 U258 ( .A(\u_div/PartRem[15][3] ), .B(\u_div/PartRem[15][2] ), .Y(
        \u_div/SumTmp[14][3] ) );
  OR2X1 U259 ( .A(\u_div/PartRem[15][2] ), .B(\u_div/PartRem[15][3] ), .Y(
        \u_div/u_add_PartRem_2_14/n3 ) );
  OR2X1 U260 ( .A(\u_div/PartRem[14][5] ), .B(\u_div/u_add_PartRem_2_13/n2 ), 
        .Y(\u_div/CryTmp[13][6] ) );
  OR2X1 U261 ( .A(\u_div/PartRem[13][5] ), .B(\u_div/u_add_PartRem_2_12/n2 ), 
        .Y(\u_div/CryTmp[12][6] ) );
  OR2X1 U262 ( .A(\u_div/PartRem[12][5] ), .B(\u_div/u_add_PartRem_2_11/n2 ), 
        .Y(\u_div/CryTmp[11][6] ) );
  OR2X1 U263 ( .A(\u_div/PartRem[11][5] ), .B(\u_div/u_add_PartRem_2_10/n2 ), 
        .Y(\u_div/CryTmp[10][6] ) );
  OR2X1 U264 ( .A(\u_div/PartRem[10][5] ), .B(\u_div/u_add_PartRem_2_9/n2 ), 
        .Y(\u_div/CryTmp[9][6] ) );
  OR2X1 U265 ( .A(\u_div/PartRem[9][5] ), .B(\u_div/u_add_PartRem_2_8/n2 ), 
        .Y(\u_div/CryTmp[8][6] ) );
  OR2X1 U266 ( .A(\u_div/PartRem[8][5] ), .B(\u_div/u_add_PartRem_2_7/n2 ), 
        .Y(\u_div/CryTmp[7][6] ) );
  OR2X1 U267 ( .A(\u_div/PartRem[7][5] ), .B(\u_div/u_add_PartRem_2_6/n2 ), 
        .Y(\u_div/CryTmp[6][6] ) );
  OR2X1 U268 ( .A(\u_div/PartRem[6][5] ), .B(\u_div/u_add_PartRem_2_5/n2 ), 
        .Y(\u_div/CryTmp[5][6] ) );
  OR2X1 U269 ( .A(\u_div/PartRem[5][5] ), .B(\u_div/u_add_PartRem_2_4/n2 ), 
        .Y(\u_div/CryTmp[4][6] ) );
  OR2X1 U270 ( .A(\u_div/PartRem[4][5] ), .B(\u_div/u_add_PartRem_2_3/n2 ), 
        .Y(\u_div/CryTmp[3][6] ) );
  OR2X1 U271 ( .A(\u_div/PartRem[3][5] ), .B(\u_div/u_add_PartRem_2_2/n2 ), 
        .Y(\u_div/CryTmp[2][6] ) );
  OR2X1 U272 ( .A(\u_div/PartRem[2][5] ), .B(\u_div/u_add_PartRem_2_1/n2 ), 
        .Y(\u_div/CryTmp[1][6] ) );
  AO21X1 U273 ( .A0(\u_div/PartRem[1][4] ), .A1(\u_div/CryTmp[1][6] ), .B0(
        \u_div/PartRem[1][5] ), .Y(\u_div/CryTmp[0][6] ) );
  NOR2X1 U274 ( .A(\u_div/PartRem[63][0] ), .B(\u_div/PartRem[62][0] ), .Y(n6)
         );
  XNOR2X1 U275 ( .A(\u_div/PartRem[63][0] ), .B(\u_div/PartRem[62][0] ), .Y(
        \u_div/SumTmp[59][3] ) );
  XNOR2X1 U276 ( .A(\u_div/PartRem[64][0] ), .B(n6), .Y(\u_div/SumTmp[59][4] )
         );
  XOR2X1 U277 ( .A(\u_div/CryTmp[9][6] ), .B(n2), .Y(\u_div/QInv[9] ) );
  XOR2X1 U278 ( .A(\u_div/CryTmp[8][6] ), .B(n3), .Y(\u_div/QInv[8] ) );
  XOR2X1 U279 ( .A(\u_div/CryTmp[7][6] ), .B(n2), .Y(\u_div/QInv[7] ) );
  XOR2X1 U280 ( .A(\u_div/CryTmp[6][6] ), .B(n3), .Y(\u_div/QInv[6] ) );
  XOR2X1 U281 ( .A(\u_div/CryTmp[5][6] ), .B(n3), .Y(\u_div/QInv[5] ) );
  XOR2X1 U282 ( .A(\u_div/CryTmp[58][6] ), .B(n3), .Y(\u_div/QInv[58] ) );
  XOR2X1 U283 ( .A(\u_div/CryTmp[57][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[57] ) );
  XOR2X1 U284 ( .A(\u_div/CryTmp[56][6] ), .B(n2), .Y(\u_div/QInv[56] ) );
  XOR2X1 U285 ( .A(\u_div/CryTmp[55][6] ), .B(n3), .Y(\u_div/QInv[55] ) );
  XOR2X1 U286 ( .A(\u_div/CryTmp[54][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[54] ) );
  XOR2X1 U287 ( .A(\u_div/CryTmp[53][6] ), .B(n2), .Y(\u_div/QInv[53] ) );
  XOR2X1 U288 ( .A(\u_div/CryTmp[52][6] ), .B(n3), .Y(\u_div/QInv[52] ) );
  XOR2X1 U289 ( .A(\u_div/CryTmp[51][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[51] ) );
  XOR2X1 U290 ( .A(\u_div/CryTmp[50][6] ), .B(n2), .Y(\u_div/QInv[50] ) );
  XOR2X1 U291 ( .A(\u_div/CryTmp[4][6] ), .B(n3), .Y(\u_div/QInv[4] ) );
  XOR2X1 U292 ( .A(\u_div/CryTmp[49][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[49] ) );
  XOR2X1 U293 ( .A(\u_div/CryTmp[48][6] ), .B(n2), .Y(\u_div/QInv[48] ) );
  XOR2X1 U294 ( .A(\u_div/CryTmp[47][6] ), .B(n3), .Y(\u_div/QInv[47] ) );
  XOR2X1 U295 ( .A(\u_div/CryTmp[46][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[46] ) );
  XOR2X1 U296 ( .A(\u_div/CryTmp[45][6] ), .B(n2), .Y(\u_div/QInv[45] ) );
  XOR2X1 U297 ( .A(\u_div/CryTmp[44][6] ), .B(n3), .Y(\u_div/QInv[44] ) );
  XOR2X1 U298 ( .A(\u_div/CryTmp[43][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[43] ) );
  XOR2X1 U299 ( .A(\u_div/CryTmp[42][6] ), .B(n2), .Y(\u_div/QInv[42] ) );
  XOR2X1 U300 ( .A(\u_div/CryTmp[41][6] ), .B(n3), .Y(\u_div/QInv[41] ) );
  XOR2X1 U301 ( .A(\u_div/CryTmp[40][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[40] ) );
  XOR2X1 U302 ( .A(\u_div/CryTmp[3][6] ), .B(n2), .Y(\u_div/QInv[3] ) );
  XOR2X1 U303 ( .A(\u_div/CryTmp[39][6] ), .B(n3), .Y(\u_div/QInv[39] ) );
  XOR2X1 U304 ( .A(\u_div/CryTmp[38][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[38] ) );
  XOR2X1 U305 ( .A(\u_div/CryTmp[37][6] ), .B(n2), .Y(\u_div/QInv[37] ) );
  XOR2X1 U306 ( .A(\u_div/CryTmp[36][6] ), .B(n3), .Y(\u_div/QInv[36] ) );
  XOR2X1 U307 ( .A(\u_div/CryTmp[35][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[35] ) );
  XOR2X1 U308 ( .A(\u_div/CryTmp[34][6] ), .B(n3), .Y(\u_div/QInv[34] ) );
  XOR2X1 U309 ( .A(\u_div/CryTmp[33][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[33] ) );
  XOR2X1 U310 ( .A(\u_div/CryTmp[32][6] ), .B(n2), .Y(\u_div/QInv[32] ) );
  XOR2X1 U311 ( .A(\u_div/CryTmp[31][6] ), .B(n3), .Y(\u_div/QInv[31] ) );
  XOR2X1 U312 ( .A(\u_div/CryTmp[30][6] ), .B(\u_div/QInv[63] ), .Y(
        \u_div/QInv[30] ) );
  XOR2X1 U313 ( .A(\u_div/CryTmp[2][6] ), .B(n2), .Y(\u_div/QInv[2] ) );
  XOR2X1 U314 ( .A(\u_div/CryTmp[29][6] ), .B(n3), .Y(\u_div/QInv[29] ) );
  XOR2X1 U315 ( .A(\u_div/CryTmp[28][6] ), .B(n4), .Y(\u_div/QInv[28] ) );
  XOR2X1 U316 ( .A(\u_div/CryTmp[27][6] ), .B(n2), .Y(\u_div/QInv[27] ) );
  XOR2X1 U317 ( .A(\u_div/CryTmp[26][6] ), .B(n3), .Y(\u_div/QInv[26] ) );
  XOR2X1 U318 ( .A(\u_div/CryTmp[25][6] ), .B(n4), .Y(\u_div/QInv[25] ) );
  XOR2X1 U319 ( .A(\u_div/CryTmp[24][6] ), .B(n2), .Y(\u_div/QInv[24] ) );
  XOR2X1 U320 ( .A(\u_div/CryTmp[23][6] ), .B(n3), .Y(\u_div/QInv[23] ) );
  XOR2X1 U321 ( .A(\u_div/CryTmp[22][6] ), .B(n4), .Y(\u_div/QInv[22] ) );
  XOR2X1 U322 ( .A(\u_div/CryTmp[21][6] ), .B(n2), .Y(\u_div/QInv[21] ) );
  XOR2X1 U323 ( .A(\u_div/CryTmp[20][6] ), .B(n3), .Y(\u_div/QInv[20] ) );
  XOR2X1 U324 ( .A(\u_div/CryTmp[1][6] ), .B(n3), .Y(\u_div/QInv[1] ) );
  XOR2X1 U325 ( .A(\u_div/CryTmp[19][6] ), .B(n2), .Y(\u_div/QInv[19] ) );
  XOR2X1 U326 ( .A(\u_div/CryTmp[18][6] ), .B(n3), .Y(\u_div/QInv[18] ) );
  XOR2X1 U327 ( .A(\u_div/CryTmp[17][6] ), .B(n4), .Y(\u_div/QInv[17] ) );
  XOR2X1 U328 ( .A(\u_div/CryTmp[16][6] ), .B(n3), .Y(\u_div/QInv[16] ) );
  XOR2X1 U329 ( .A(\u_div/CryTmp[15][6] ), .B(n4), .Y(\u_div/QInv[15] ) );
  XOR2X1 U330 ( .A(\u_div/CryTmp[14][6] ), .B(n3), .Y(\u_div/QInv[14] ) );
  XOR2X1 U331 ( .A(\u_div/CryTmp[13][6] ), .B(n4), .Y(\u_div/QInv[13] ) );
  XOR2X1 U332 ( .A(\u_div/CryTmp[12][6] ), .B(n3), .Y(\u_div/QInv[12] ) );
  XOR2X1 U333 ( .A(\u_div/CryTmp[11][6] ), .B(n2), .Y(\u_div/QInv[11] ) );
  XOR2X1 U334 ( .A(\u_div/CryTmp[10][6] ), .B(n3), .Y(\u_div/QInv[10] ) );
  XOR2X1 U335 ( .A(\u_div/CryTmp[0][6] ), .B(n3), .Y(\u_div/QInv[0] ) );
endmodule


module GSIM_DW01_inc_10 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  ADDHXL U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  ADDHXL U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  ADDHXL U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  ADDHXL U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  ADDHXL U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  ADDHXL U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  ADDHXL U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  ADDHXL U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  ADDHXL U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  ADDHXL U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  ADDHXL U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  ADDHXL U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[31]), .B(A[31]), .Y(SUM[31]) );
endmodule


module GSIM_DW01_inc_11 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  ADDHXL U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  ADDHX1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHX1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHX1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHX1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHX1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  ADDHXL U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  ADDHXL U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  ADDHXL U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  ADDHXL U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  ADDHXL U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[31]), .B(A[31]), .Y(SUM[31]) );
endmodule


module GSIM_DW_mult_tc_21 ( a, b, product );
  input [4:0] a;
  input [63:0] b;
  output [68:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, \b[0] , \b[1] , n321, n322, n323;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[1] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U3 ( .A(n65), .B(n66), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U4 ( .A(n67), .B(n68), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U14 ( .A(n87), .B(n88), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U16 ( .A(n91), .B(n92), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U18 ( .A(n95), .B(n96), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U20 ( .A(n99), .B(n100), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U22 ( .A(n103), .B(n104), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U24 ( .A(n107), .B(n108), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U26 ( .A(n111), .B(n112), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U28 ( .A(n115), .B(n116), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U30 ( .A(n119), .B(n120), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U50 ( .A(n159), .B(n160), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U52 ( .A(n163), .B(n164), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U54 ( .A(n167), .B(n168), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U56 ( .A(n171), .B(n172), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U58 ( .A(n175), .B(n176), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U60 ( .A(n179), .B(n180), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U62 ( .A(n62), .B(\b[0] ), .CI(n183), .CO(n61), .S(product[3]) );
  ADDHXL U63 ( .A(\b[0] ), .B(b[2]), .CO(n62), .S(product[2]) );
  ADDFXL U65 ( .A(b[59]), .B(b[62]), .CI(b[60]), .CO(n64), .S(n65) );
  ADDFXL U66 ( .A(b[58]), .B(b[61]), .CI(b[59]), .CO(n66), .S(n67) );
  ADDFXL U67 ( .A(b[57]), .B(b[60]), .CI(b[58]), .CO(n68), .S(n69) );
  ADDFXL U68 ( .A(b[56]), .B(b[59]), .CI(b[57]), .CO(n70), .S(n71) );
  ADDFXL U69 ( .A(b[55]), .B(b[58]), .CI(b[56]), .CO(n72), .S(n73) );
  ADDFXL U70 ( .A(b[54]), .B(b[57]), .CI(b[55]), .CO(n74), .S(n75) );
  ADDFXL U71 ( .A(b[53]), .B(b[56]), .CI(b[54]), .CO(n76), .S(n77) );
  ADDFXL U72 ( .A(b[52]), .B(b[55]), .CI(b[53]), .CO(n78), .S(n79) );
  ADDFXL U73 ( .A(b[51]), .B(b[54]), .CI(b[52]), .CO(n80), .S(n81) );
  ADDFXL U74 ( .A(b[50]), .B(b[53]), .CI(b[51]), .CO(n82), .S(n83) );
  ADDFXL U75 ( .A(b[49]), .B(b[52]), .CI(b[50]), .CO(n84), .S(n85) );
  ADDFXL U76 ( .A(b[48]), .B(b[51]), .CI(b[49]), .CO(n86), .S(n87) );
  ADDFXL U77 ( .A(b[47]), .B(b[50]), .CI(b[48]), .CO(n88), .S(n89) );
  ADDFXL U78 ( .A(b[46]), .B(b[49]), .CI(b[47]), .CO(n90), .S(n91) );
  ADDFXL U79 ( .A(b[45]), .B(b[48]), .CI(b[46]), .CO(n92), .S(n93) );
  ADDFXL U80 ( .A(b[44]), .B(b[47]), .CI(b[45]), .CO(n94), .S(n95) );
  ADDFXL U81 ( .A(b[43]), .B(b[46]), .CI(b[44]), .CO(n96), .S(n97) );
  ADDFXL U82 ( .A(b[42]), .B(b[45]), .CI(b[43]), .CO(n98), .S(n99) );
  ADDFXL U83 ( .A(b[41]), .B(b[44]), .CI(b[42]), .CO(n100), .S(n101) );
  ADDFXL U84 ( .A(b[40]), .B(b[43]), .CI(b[41]), .CO(n102), .S(n103) );
  ADDFXL U85 ( .A(b[39]), .B(b[42]), .CI(b[40]), .CO(n104), .S(n105) );
  ADDFXL U86 ( .A(b[38]), .B(b[41]), .CI(b[39]), .CO(n106), .S(n107) );
  ADDFXL U87 ( .A(b[37]), .B(b[40]), .CI(b[38]), .CO(n108), .S(n109) );
  ADDFXL U88 ( .A(b[36]), .B(b[39]), .CI(b[37]), .CO(n110), .S(n111) );
  ADDFXL U89 ( .A(b[35]), .B(b[38]), .CI(b[36]), .CO(n112), .S(n113) );
  ADDFXL U90 ( .A(b[34]), .B(b[37]), .CI(b[35]), .CO(n114), .S(n115) );
  ADDFXL U91 ( .A(b[33]), .B(b[36]), .CI(b[34]), .CO(n116), .S(n117) );
  ADDFXL U92 ( .A(b[32]), .B(b[35]), .CI(b[33]), .CO(n118), .S(n119) );
  ADDFXL U93 ( .A(b[31]), .B(b[34]), .CI(b[32]), .CO(n120), .S(n121) );
  ADDFXL U94 ( .A(b[30]), .B(b[33]), .CI(b[31]), .CO(n122), .S(n123) );
  ADDFXL U95 ( .A(b[29]), .B(b[32]), .CI(b[30]), .CO(n124), .S(n125) );
  ADDFXL U96 ( .A(b[28]), .B(b[31]), .CI(b[29]), .CO(n126), .S(n127) );
  ADDFXL U97 ( .A(b[27]), .B(b[30]), .CI(b[28]), .CO(n128), .S(n129) );
  ADDFXL U98 ( .A(b[26]), .B(b[29]), .CI(b[27]), .CO(n130), .S(n131) );
  ADDFXL U99 ( .A(b[25]), .B(b[28]), .CI(b[26]), .CO(n132), .S(n133) );
  ADDFXL U100 ( .A(b[24]), .B(b[27]), .CI(b[25]), .CO(n134), .S(n135) );
  ADDFXL U101 ( .A(b[23]), .B(b[26]), .CI(b[24]), .CO(n136), .S(n137) );
  ADDFXL U102 ( .A(b[22]), .B(b[25]), .CI(b[23]), .CO(n138), .S(n139) );
  ADDFXL U103 ( .A(b[21]), .B(b[24]), .CI(b[22]), .CO(n140), .S(n141) );
  ADDFXL U104 ( .A(b[20]), .B(b[23]), .CI(b[21]), .CO(n142), .S(n143) );
  ADDFXL U105 ( .A(b[19]), .B(b[22]), .CI(b[20]), .CO(n144), .S(n145) );
  ADDFXL U106 ( .A(b[18]), .B(b[21]), .CI(b[19]), .CO(n146), .S(n147) );
  ADDFXL U107 ( .A(b[17]), .B(b[20]), .CI(b[18]), .CO(n148), .S(n149) );
  ADDFXL U108 ( .A(b[16]), .B(b[19]), .CI(b[17]), .CO(n150), .S(n151) );
  ADDFXL U109 ( .A(b[15]), .B(b[18]), .CI(b[16]), .CO(n152), .S(n153) );
  ADDFXL U110 ( .A(b[14]), .B(b[17]), .CI(b[15]), .CO(n154), .S(n155) );
  ADDFXL U111 ( .A(b[13]), .B(b[16]), .CI(b[14]), .CO(n156), .S(n157) );
  ADDFXL U112 ( .A(b[12]), .B(b[15]), .CI(b[13]), .CO(n158), .S(n159) );
  ADDFXL U113 ( .A(b[11]), .B(b[14]), .CI(b[12]), .CO(n160), .S(n161) );
  ADDFXL U114 ( .A(b[10]), .B(b[13]), .CI(b[11]), .CO(n162), .S(n163) );
  ADDFXL U115 ( .A(b[9]), .B(b[12]), .CI(b[10]), .CO(n164), .S(n165) );
  ADDFXL U116 ( .A(b[8]), .B(b[11]), .CI(b[9]), .CO(n166), .S(n167) );
  ADDFXL U117 ( .A(b[7]), .B(b[10]), .CI(b[8]), .CO(n168), .S(n169) );
  ADDFXL U118 ( .A(b[6]), .B(b[9]), .CI(b[7]), .CO(n170), .S(n171) );
  ADDFXL U119 ( .A(b[5]), .B(b[8]), .CI(b[6]), .CO(n172), .S(n173) );
  ADDFXL U120 ( .A(b[4]), .B(b[7]), .CI(b[5]), .CO(n174), .S(n175) );
  ADDFXL U121 ( .A(b[3]), .B(b[6]), .CI(b[4]), .CO(n176), .S(n177) );
  ADDFXL U122 ( .A(b[2]), .B(b[5]), .CI(b[3]), .CO(n178), .S(n179) );
  ADDHXL U124 ( .A(b[3]), .B(\b[1] ), .CO(n182), .S(n183) );
  ADDFXL U129 ( .A(n161), .B(n162), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U130 ( .A(n157), .B(n158), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U131 ( .A(n155), .B(n156), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U132 ( .A(n153), .B(n154), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U133 ( .A(n151), .B(n152), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U134 ( .A(n149), .B(n150), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U135 ( .A(n147), .B(n148), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U136 ( .A(n139), .B(n140), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U137 ( .A(n141), .B(n142), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U138 ( .A(n143), .B(n144), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U139 ( .A(n145), .B(n146), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U140 ( .A(\b[1] ), .B(b[4]), .CI(b[2]), .CO(n180), .S(n181) );
  ADDFXL U141 ( .A(n165), .B(n166), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U142 ( .A(n169), .B(n170), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U143 ( .A(n173), .B(n174), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U144 ( .A(n177), .B(n178), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U145 ( .A(n135), .B(n136), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U146 ( .A(n131), .B(n132), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U147 ( .A(n127), .B(n128), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U148 ( .A(n121), .B(n122), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U149 ( .A(n117), .B(n118), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U150 ( .A(n113), .B(n114), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U151 ( .A(n109), .B(n110), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U152 ( .A(n105), .B(n106), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U153 ( .A(n101), .B(n102), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U154 ( .A(n97), .B(n98), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U155 ( .A(n93), .B(n94), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U156 ( .A(n89), .B(n90), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U157 ( .A(n85), .B(n86), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U158 ( .A(n83), .B(n84), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U159 ( .A(n79), .B(n80), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U160 ( .A(n75), .B(n76), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U161 ( .A(n71), .B(n72), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U162 ( .A(n69), .B(n70), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U163 ( .A(n137), .B(n138), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U164 ( .A(n123), .B(n124), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U165 ( .A(n81), .B(n82), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U166 ( .A(n125), .B(n126), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U167 ( .A(n181), .B(n182), .CI(n61), .CO(n60), .S(product[4]) );
  ADDFXL U168 ( .A(n133), .B(n134), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U169 ( .A(n129), .B(n130), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U170 ( .A(n77), .B(n78), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U171 ( .A(n73), .B(n74), .CI(n7), .CO(n6), .S(product[58]) );
  XNOR2XL U172 ( .A(b[61]), .B(b[60]), .Y(n322) );
  XOR2X1 U173 ( .A(n321), .B(n322), .Y(product[63]) );
  XOR2X1 U174 ( .A(n323), .B(b[63]), .Y(n321) );
  XNOR2X1 U175 ( .A(n64), .B(n2), .Y(n323) );
endmodule


module GSIM_DW_mult_tc_20 ( a, b, product );
  input [3:0] a;
  input [63:0] b;
  output [67:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, \b[0] , \b[1] , n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318;
  assign product[1] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[2] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U3 ( .A(b[61]), .B(n317), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U4 ( .A(b[60]), .B(n316), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U5 ( .A(b[59]), .B(n315), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U6 ( .A(b[58]), .B(n314), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U7 ( .A(b[57]), .B(n313), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U8 ( .A(b[56]), .B(n312), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U9 ( .A(b[55]), .B(n311), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U10 ( .A(b[54]), .B(n310), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U11 ( .A(b[53]), .B(n309), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U12 ( .A(b[52]), .B(n308), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U13 ( .A(b[51]), .B(n307), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U14 ( .A(b[50]), .B(n306), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U15 ( .A(b[49]), .B(n305), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U16 ( .A(b[48]), .B(n304), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U17 ( .A(b[47]), .B(n303), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U18 ( .A(b[46]), .B(n302), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U19 ( .A(b[45]), .B(n301), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U20 ( .A(b[44]), .B(n300), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U21 ( .A(b[43]), .B(n299), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U22 ( .A(b[42]), .B(n298), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U23 ( .A(b[41]), .B(n297), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U24 ( .A(b[40]), .B(n296), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U25 ( .A(b[39]), .B(n295), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U26 ( .A(b[38]), .B(n294), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U27 ( .A(b[37]), .B(n293), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U28 ( .A(b[36]), .B(n292), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U29 ( .A(b[35]), .B(n291), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U30 ( .A(b[34]), .B(n290), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U31 ( .A(b[33]), .B(n289), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U32 ( .A(b[32]), .B(n288), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U33 ( .A(b[31]), .B(n287), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U34 ( .A(b[30]), .B(n286), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U35 ( .A(b[29]), .B(n285), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U36 ( .A(b[28]), .B(n284), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U37 ( .A(b[27]), .B(n283), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U38 ( .A(b[26]), .B(n282), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U39 ( .A(b[25]), .B(n281), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U40 ( .A(b[24]), .B(n280), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U41 ( .A(b[23]), .B(n279), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U42 ( .A(b[22]), .B(n278), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U43 ( .A(b[21]), .B(n277), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U44 ( .A(b[20]), .B(n276), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U45 ( .A(b[19]), .B(n275), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U46 ( .A(b[18]), .B(n274), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U47 ( .A(b[17]), .B(n273), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U48 ( .A(b[16]), .B(n272), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U49 ( .A(b[15]), .B(n271), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U50 ( .A(b[14]), .B(n270), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U51 ( .A(b[13]), .B(n269), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U52 ( .A(b[12]), .B(n268), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U53 ( .A(b[11]), .B(n267), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U54 ( .A(b[10]), .B(n266), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U55 ( .A(b[9]), .B(n265), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U56 ( .A(b[8]), .B(n264), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U57 ( .A(b[7]), .B(n263), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U58 ( .A(b[6]), .B(n262), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U59 ( .A(b[5]), .B(n261), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U60 ( .A(b[4]), .B(n260), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U61 ( .A(b[3]), .B(n259), .CI(n61), .CO(n60), .S(product[4]) );
  INVXL U131 ( .A(\b[1] ), .Y(n259) );
  INVXL U132 ( .A(b[18]), .Y(n276) );
  INVXL U133 ( .A(b[28]), .Y(n286) );
  INVXL U134 ( .A(b[38]), .Y(n296) );
  INVXL U135 ( .A(b[48]), .Y(n306) );
  INVXL U136 ( .A(b[10]), .Y(n268) );
  INVXL U137 ( .A(b[17]), .Y(n275) );
  INVXL U138 ( .A(b[19]), .Y(n277) );
  INVXL U139 ( .A(b[20]), .Y(n278) );
  INVXL U140 ( .A(b[27]), .Y(n285) );
  INVXL U141 ( .A(b[29]), .Y(n287) );
  INVXL U142 ( .A(b[30]), .Y(n288) );
  INVXL U143 ( .A(b[37]), .Y(n295) );
  INVXL U144 ( .A(b[39]), .Y(n297) );
  INVXL U145 ( .A(b[40]), .Y(n298) );
  INVXL U146 ( .A(b[47]), .Y(n305) );
  INVXL U147 ( .A(b[49]), .Y(n307) );
  INVXL U148 ( .A(b[50]), .Y(n308) );
  INVXL U149 ( .A(b[51]), .Y(n309) );
  INVXL U150 ( .A(b[6]), .Y(n264) );
  INVXL U151 ( .A(b[7]), .Y(n265) );
  INVXL U152 ( .A(b[8]), .Y(n266) );
  INVXL U153 ( .A(b[9]), .Y(n267) );
  INVXL U154 ( .A(b[16]), .Y(n274) );
  INVXL U155 ( .A(b[26]), .Y(n284) );
  INVXL U156 ( .A(b[36]), .Y(n294) );
  INVXL U157 ( .A(b[46]), .Y(n304) );
  INVXL U158 ( .A(b[3]), .Y(n261) );
  INVXL U159 ( .A(b[4]), .Y(n262) );
  INVXL U160 ( .A(b[5]), .Y(n263) );
  INVXL U161 ( .A(b[11]), .Y(n269) );
  INVXL U162 ( .A(b[12]), .Y(n270) );
  INVXL U163 ( .A(b[13]), .Y(n271) );
  INVXL U164 ( .A(b[14]), .Y(n272) );
  INVXL U165 ( .A(b[15]), .Y(n273) );
  INVXL U166 ( .A(b[21]), .Y(n279) );
  INVXL U167 ( .A(b[22]), .Y(n280) );
  INVXL U168 ( .A(b[23]), .Y(n281) );
  INVXL U169 ( .A(b[24]), .Y(n282) );
  INVXL U170 ( .A(b[25]), .Y(n283) );
  INVXL U171 ( .A(b[31]), .Y(n289) );
  INVXL U172 ( .A(b[32]), .Y(n290) );
  INVXL U173 ( .A(b[33]), .Y(n291) );
  INVXL U174 ( .A(b[34]), .Y(n292) );
  INVXL U175 ( .A(b[35]), .Y(n293) );
  INVXL U176 ( .A(b[41]), .Y(n299) );
  INVXL U177 ( .A(b[42]), .Y(n300) );
  INVXL U178 ( .A(b[43]), .Y(n301) );
  INVXL U179 ( .A(b[44]), .Y(n302) );
  INVXL U180 ( .A(b[45]), .Y(n303) );
  INVXL U181 ( .A(b[52]), .Y(n310) );
  INVXL U182 ( .A(b[53]), .Y(n311) );
  INVXL U183 ( .A(b[54]), .Y(n312) );
  INVXL U184 ( .A(b[55]), .Y(n313) );
  INVXL U185 ( .A(b[56]), .Y(n314) );
  INVXL U186 ( .A(b[57]), .Y(n315) );
  INVXL U187 ( .A(b[58]), .Y(n316) );
  INVXL U188 ( .A(b[59]), .Y(n317) );
  INVXL U189 ( .A(b[2]), .Y(n260) );
  XOR2X1 U190 ( .A(n318), .B(b[60]), .Y(product[63]) );
  XNOR2X1 U191 ( .A(n2), .B(b[62]), .Y(n318) );
  XOR2X1 U192 ( .A(b[2]), .B(\b[0] ), .Y(product[3]) );
  NAND2X1 U193 ( .A(\b[0] ), .B(n260), .Y(n61) );
endmodule


module GSIM_DW_mult_tc_19 ( a, b, product );
  input [3:0] a;
  input [63:0] b;
  output [67:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, \b[0] , \b[1] , n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318;
  assign product[1] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[2] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U3 ( .A(b[61]), .B(n317), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U4 ( .A(b[60]), .B(n316), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U5 ( .A(b[59]), .B(n315), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U6 ( .A(b[58]), .B(n314), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U7 ( .A(b[57]), .B(n313), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U8 ( .A(b[56]), .B(n312), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U9 ( .A(b[55]), .B(n311), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U10 ( .A(b[54]), .B(n310), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U11 ( .A(b[53]), .B(n309), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U12 ( .A(b[52]), .B(n308), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U13 ( .A(b[51]), .B(n307), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U14 ( .A(b[50]), .B(n306), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U15 ( .A(b[49]), .B(n305), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U16 ( .A(b[48]), .B(n304), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U17 ( .A(b[47]), .B(n303), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U18 ( .A(b[46]), .B(n302), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U19 ( .A(b[45]), .B(n301), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U20 ( .A(b[44]), .B(n300), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U21 ( .A(b[43]), .B(n299), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U22 ( .A(b[42]), .B(n298), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U23 ( .A(b[41]), .B(n297), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U24 ( .A(b[40]), .B(n296), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U25 ( .A(b[39]), .B(n295), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U26 ( .A(b[38]), .B(n294), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U27 ( .A(b[37]), .B(n293), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U28 ( .A(b[36]), .B(n292), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U29 ( .A(b[35]), .B(n291), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U30 ( .A(b[34]), .B(n290), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U31 ( .A(b[33]), .B(n289), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U32 ( .A(b[32]), .B(n288), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U33 ( .A(b[31]), .B(n287), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U34 ( .A(b[30]), .B(n286), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U35 ( .A(b[29]), .B(n285), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U36 ( .A(b[28]), .B(n284), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U37 ( .A(b[27]), .B(n283), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U38 ( .A(b[26]), .B(n282), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U39 ( .A(b[25]), .B(n281), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U40 ( .A(b[24]), .B(n280), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U41 ( .A(b[23]), .B(n279), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U42 ( .A(b[22]), .B(n278), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U43 ( .A(b[21]), .B(n277), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U44 ( .A(b[20]), .B(n276), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U45 ( .A(b[19]), .B(n275), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U46 ( .A(b[18]), .B(n274), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U47 ( .A(b[17]), .B(n273), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U48 ( .A(b[16]), .B(n272), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U49 ( .A(b[15]), .B(n271), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U50 ( .A(b[14]), .B(n270), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U51 ( .A(b[13]), .B(n269), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U52 ( .A(b[12]), .B(n268), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U53 ( .A(b[11]), .B(n267), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U54 ( .A(b[10]), .B(n266), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U55 ( .A(b[9]), .B(n265), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U56 ( .A(b[8]), .B(n264), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U57 ( .A(b[7]), .B(n263), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U58 ( .A(b[6]), .B(n262), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U59 ( .A(b[5]), .B(n261), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U60 ( .A(b[4]), .B(n260), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U61 ( .A(b[3]), .B(n259), .CI(n61), .CO(n60), .S(product[4]) );
  CLKINVX1 U131 ( .A(\b[1] ), .Y(n259) );
  NAND2X1 U132 ( .A(\b[0] ), .B(n260), .Y(n61) );
  INVXL U133 ( .A(b[2]), .Y(n260) );
  XOR2XL U134 ( .A(b[2]), .B(\b[0] ), .Y(product[3]) );
  INVXL U135 ( .A(b[42]), .Y(n300) );
  INVXL U136 ( .A(b[41]), .Y(n299) );
  INVXL U137 ( .A(b[32]), .Y(n290) );
  INVXL U138 ( .A(b[31]), .Y(n289) );
  INVXL U139 ( .A(b[21]), .Y(n279) );
  INVXL U140 ( .A(b[22]), .Y(n280) );
  INVXL U141 ( .A(b[12]), .Y(n270) );
  INVXL U142 ( .A(b[11]), .Y(n269) );
  CLKINVX1 U143 ( .A(b[52]), .Y(n310) );
  INVXL U144 ( .A(b[4]), .Y(n262) );
  INVXL U145 ( .A(b[3]), .Y(n261) );
  CLKINVX1 U146 ( .A(b[51]), .Y(n309) );
  INVXL U147 ( .A(b[14]), .Y(n272) );
  INVXL U148 ( .A(b[24]), .Y(n282) );
  INVXL U149 ( .A(b[34]), .Y(n292) );
  INVXL U150 ( .A(b[44]), .Y(n302) );
  INVXL U151 ( .A(b[54]), .Y(n312) );
  INVXL U152 ( .A(b[5]), .Y(n263) );
  INVXL U153 ( .A(b[6]), .Y(n264) );
  INVXL U154 ( .A(b[7]), .Y(n265) );
  INVXL U155 ( .A(b[8]), .Y(n266) );
  INVXL U156 ( .A(b[9]), .Y(n267) );
  INVXL U157 ( .A(b[10]), .Y(n268) );
  INVXL U158 ( .A(b[13]), .Y(n271) );
  INVXL U159 ( .A(b[15]), .Y(n273) );
  INVXL U160 ( .A(b[16]), .Y(n274) );
  INVXL U161 ( .A(b[17]), .Y(n275) );
  INVXL U162 ( .A(b[18]), .Y(n276) );
  INVXL U163 ( .A(b[19]), .Y(n277) );
  INVXL U164 ( .A(b[20]), .Y(n278) );
  INVXL U165 ( .A(b[23]), .Y(n281) );
  INVXL U166 ( .A(b[25]), .Y(n283) );
  INVXL U167 ( .A(b[26]), .Y(n284) );
  INVXL U168 ( .A(b[27]), .Y(n285) );
  INVXL U169 ( .A(b[28]), .Y(n286) );
  INVXL U170 ( .A(b[29]), .Y(n287) );
  INVXL U171 ( .A(b[30]), .Y(n288) );
  INVXL U172 ( .A(b[33]), .Y(n291) );
  INVXL U173 ( .A(b[35]), .Y(n293) );
  INVXL U174 ( .A(b[36]), .Y(n294) );
  INVXL U175 ( .A(b[37]), .Y(n295) );
  INVXL U176 ( .A(b[38]), .Y(n296) );
  INVXL U177 ( .A(b[39]), .Y(n297) );
  INVXL U178 ( .A(b[40]), .Y(n298) );
  INVXL U179 ( .A(b[43]), .Y(n301) );
  INVXL U180 ( .A(b[45]), .Y(n303) );
  INVXL U181 ( .A(b[46]), .Y(n304) );
  INVXL U182 ( .A(b[47]), .Y(n305) );
  INVXL U183 ( .A(b[48]), .Y(n306) );
  INVXL U184 ( .A(b[49]), .Y(n307) );
  INVXL U185 ( .A(b[50]), .Y(n308) );
  INVXL U186 ( .A(b[53]), .Y(n311) );
  INVXL U187 ( .A(b[55]), .Y(n313) );
  INVXL U188 ( .A(b[56]), .Y(n314) );
  INVXL U189 ( .A(b[57]), .Y(n315) );
  INVXL U190 ( .A(b[58]), .Y(n316) );
  CLKINVX1 U191 ( .A(b[59]), .Y(n317) );
  XOR2X1 U192 ( .A(n318), .B(b[60]), .Y(product[63]) );
  XNOR2X1 U193 ( .A(n2), .B(b[62]), .Y(n318) );
endmodule


module GSIM_DW01_add_501 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;
  assign SUM[15] = B[15];
  assign SUM[14] = B[14];
  assign SUM[13] = B[13];
  assign SUM[12] = B[12];
  assign SUM[11] = B[11];
  assign SUM[10] = B[10];
  assign SUM[9] = B[9];
  assign SUM[8] = B[8];
  assign SUM[7] = B[7];
  assign SUM[6] = B[6];
  assign SUM[5] = B[5];
  assign SUM[4] = B[4];
  assign SUM[3] = B[3];
  assign SUM[2] = B[2];
  assign SUM[1] = B[1];

  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(n1), .CO(carry[18]), .S(SUM[17]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  AND2X2 U1 ( .A(B[16]), .B(A[16]), .Y(n1) );
  XOR2XL U2 ( .A(B[16]), .B(A[16]), .Y(SUM[16]) );
endmodule


module GSIM_DW01_add_500 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;

  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2XL U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module GSIM_DW_mult_tc_18 ( a, b, product );
  input [4:0] a;
  input [63:0] b;
  output [68:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, \b[0] , \b[1] , n321, n322, n323;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[1] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U4 ( .A(n67), .B(n68), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U7 ( .A(n73), .B(n74), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U13 ( .A(n85), .B(n86), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U15 ( .A(n89), .B(n90), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U17 ( .A(n93), .B(n94), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U19 ( .A(n97), .B(n98), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U21 ( .A(n101), .B(n102), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U23 ( .A(n105), .B(n106), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U25 ( .A(n109), .B(n110), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U27 ( .A(n113), .B(n114), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U29 ( .A(n117), .B(n118), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U49 ( .A(n157), .B(n158), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U51 ( .A(n161), .B(n162), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U53 ( .A(n165), .B(n166), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U55 ( .A(n169), .B(n170), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U57 ( .A(n173), .B(n174), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U59 ( .A(n177), .B(n178), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U61 ( .A(n181), .B(n182), .CI(n61), .CO(n60), .S(product[4]) );
  ADDHXL U63 ( .A(\b[0] ), .B(b[2]), .CO(n62), .S(product[2]) );
  ADDFXL U65 ( .A(b[59]), .B(b[62]), .CI(b[60]), .CO(n64), .S(n65) );
  ADDFXL U66 ( .A(b[58]), .B(b[61]), .CI(b[59]), .CO(n66), .S(n67) );
  ADDFXL U67 ( .A(b[57]), .B(b[60]), .CI(b[58]), .CO(n68), .S(n69) );
  ADDFXL U68 ( .A(b[56]), .B(b[59]), .CI(b[57]), .CO(n70), .S(n71) );
  ADDFXL U69 ( .A(b[55]), .B(b[58]), .CI(b[56]), .CO(n72), .S(n73) );
  ADDFXL U70 ( .A(b[54]), .B(b[57]), .CI(b[55]), .CO(n74), .S(n75) );
  ADDFXL U71 ( .A(b[53]), .B(b[56]), .CI(b[54]), .CO(n76), .S(n77) );
  ADDFXL U72 ( .A(b[52]), .B(b[55]), .CI(b[53]), .CO(n78), .S(n79) );
  ADDFXL U73 ( .A(b[51]), .B(b[54]), .CI(b[52]), .CO(n80), .S(n81) );
  ADDFXL U74 ( .A(b[50]), .B(b[53]), .CI(b[51]), .CO(n82), .S(n83) );
  ADDFXL U75 ( .A(b[49]), .B(b[52]), .CI(b[50]), .CO(n84), .S(n85) );
  ADDFXL U76 ( .A(b[48]), .B(b[51]), .CI(b[49]), .CO(n86), .S(n87) );
  ADDFXL U77 ( .A(b[47]), .B(b[50]), .CI(b[48]), .CO(n88), .S(n89) );
  ADDFXL U78 ( .A(b[46]), .B(b[49]), .CI(b[47]), .CO(n90), .S(n91) );
  ADDFXL U79 ( .A(b[45]), .B(b[48]), .CI(b[46]), .CO(n92), .S(n93) );
  ADDFXL U80 ( .A(b[44]), .B(b[47]), .CI(b[45]), .CO(n94), .S(n95) );
  ADDFXL U81 ( .A(b[43]), .B(b[46]), .CI(b[44]), .CO(n96), .S(n97) );
  ADDFXL U82 ( .A(b[42]), .B(b[45]), .CI(b[43]), .CO(n98), .S(n99) );
  ADDFXL U83 ( .A(b[41]), .B(b[44]), .CI(b[42]), .CO(n100), .S(n101) );
  ADDFXL U84 ( .A(b[40]), .B(b[43]), .CI(b[41]), .CO(n102), .S(n103) );
  ADDFXL U85 ( .A(b[39]), .B(b[42]), .CI(b[40]), .CO(n104), .S(n105) );
  ADDFXL U86 ( .A(b[38]), .B(b[41]), .CI(b[39]), .CO(n106), .S(n107) );
  ADDFXL U87 ( .A(b[37]), .B(b[40]), .CI(b[38]), .CO(n108), .S(n109) );
  ADDFXL U88 ( .A(b[36]), .B(b[39]), .CI(b[37]), .CO(n110), .S(n111) );
  ADDFXL U89 ( .A(b[35]), .B(b[38]), .CI(b[36]), .CO(n112), .S(n113) );
  ADDFXL U90 ( .A(b[34]), .B(b[37]), .CI(b[35]), .CO(n114), .S(n115) );
  ADDFXL U91 ( .A(b[33]), .B(b[36]), .CI(b[34]), .CO(n116), .S(n117) );
  ADDFXL U92 ( .A(b[32]), .B(b[35]), .CI(b[33]), .CO(n118), .S(n119) );
  ADDFXL U93 ( .A(b[31]), .B(b[34]), .CI(b[32]), .CO(n120), .S(n121) );
  ADDFXL U94 ( .A(b[30]), .B(b[33]), .CI(b[31]), .CO(n122), .S(n123) );
  ADDFXL U95 ( .A(b[29]), .B(b[32]), .CI(b[30]), .CO(n124), .S(n125) );
  ADDFXL U96 ( .A(b[28]), .B(b[31]), .CI(b[29]), .CO(n126), .S(n127) );
  ADDFXL U97 ( .A(b[27]), .B(b[30]), .CI(b[28]), .CO(n128), .S(n129) );
  ADDFXL U98 ( .A(b[26]), .B(b[29]), .CI(b[27]), .CO(n130), .S(n131) );
  ADDFXL U99 ( .A(b[25]), .B(b[28]), .CI(b[26]), .CO(n132), .S(n133) );
  ADDFXL U100 ( .A(b[24]), .B(b[27]), .CI(b[25]), .CO(n134), .S(n135) );
  ADDFXL U101 ( .A(b[23]), .B(b[26]), .CI(b[24]), .CO(n136), .S(n137) );
  ADDFXL U102 ( .A(b[22]), .B(b[25]), .CI(b[23]), .CO(n138), .S(n139) );
  ADDFXL U103 ( .A(b[21]), .B(b[24]), .CI(b[22]), .CO(n140), .S(n141) );
  ADDFXL U104 ( .A(b[20]), .B(b[23]), .CI(b[21]), .CO(n142), .S(n143) );
  ADDFXL U105 ( .A(b[19]), .B(b[22]), .CI(b[20]), .CO(n144), .S(n145) );
  ADDFXL U106 ( .A(b[18]), .B(b[21]), .CI(b[19]), .CO(n146), .S(n147) );
  ADDFXL U107 ( .A(b[17]), .B(b[20]), .CI(b[18]), .CO(n148), .S(n149) );
  ADDFXL U108 ( .A(b[16]), .B(b[19]), .CI(b[17]), .CO(n150), .S(n151) );
  ADDFXL U109 ( .A(b[15]), .B(b[18]), .CI(b[16]), .CO(n152), .S(n153) );
  ADDFXL U110 ( .A(b[14]), .B(b[17]), .CI(b[15]), .CO(n154), .S(n155) );
  ADDFXL U111 ( .A(b[13]), .B(b[16]), .CI(b[14]), .CO(n156), .S(n157) );
  ADDFXL U112 ( .A(b[12]), .B(b[15]), .CI(b[13]), .CO(n158), .S(n159) );
  ADDFXL U113 ( .A(b[11]), .B(b[14]), .CI(b[12]), .CO(n160), .S(n161) );
  ADDFXL U114 ( .A(b[10]), .B(b[13]), .CI(b[11]), .CO(n162), .S(n163) );
  ADDFXL U115 ( .A(b[9]), .B(b[12]), .CI(b[10]), .CO(n164), .S(n165) );
  ADDFXL U116 ( .A(b[8]), .B(b[11]), .CI(b[9]), .CO(n166), .S(n167) );
  ADDFXL U117 ( .A(b[7]), .B(b[10]), .CI(b[8]), .CO(n168), .S(n169) );
  ADDFXL U118 ( .A(b[6]), .B(b[9]), .CI(b[7]), .CO(n170), .S(n171) );
  ADDFXL U119 ( .A(b[5]), .B(b[8]), .CI(b[6]), .CO(n172), .S(n173) );
  ADDFXL U120 ( .A(b[4]), .B(b[7]), .CI(b[5]), .CO(n174), .S(n175) );
  ADDFXL U121 ( .A(b[3]), .B(b[6]), .CI(b[4]), .CO(n176), .S(n177) );
  ADDFXL U122 ( .A(b[2]), .B(b[5]), .CI(b[3]), .CO(n178), .S(n179) );
  ADDFXL U123 ( .A(\b[1] ), .B(b[4]), .CI(b[2]), .CO(n180), .S(n181) );
  ADDHXL U124 ( .A(b[3]), .B(\b[1] ), .CO(n182), .S(n183) );
  ADDFXL U129 ( .A(n159), .B(n160), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U130 ( .A(n155), .B(n156), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U131 ( .A(n153), .B(n154), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U132 ( .A(n151), .B(n152), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U133 ( .A(n149), .B(n150), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U134 ( .A(n147), .B(n148), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U135 ( .A(n139), .B(n140), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U136 ( .A(n141), .B(n142), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U137 ( .A(n143), .B(n144), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U138 ( .A(n145), .B(n146), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U139 ( .A(n163), .B(n164), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U140 ( .A(n179), .B(n180), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U141 ( .A(n171), .B(n172), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U142 ( .A(n167), .B(n168), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U143 ( .A(n175), .B(n176), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U144 ( .A(n137), .B(n138), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U145 ( .A(n135), .B(n136), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U146 ( .A(n133), .B(n134), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U147 ( .A(n131), .B(n132), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U148 ( .A(n129), .B(n130), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U149 ( .A(n127), .B(n128), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U150 ( .A(n125), .B(n126), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U151 ( .A(n123), .B(n124), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U152 ( .A(n119), .B(n120), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U153 ( .A(n115), .B(n116), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U154 ( .A(n111), .B(n112), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U155 ( .A(n107), .B(n108), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U156 ( .A(n103), .B(n104), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U157 ( .A(n99), .B(n100), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U158 ( .A(n95), .B(n96), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U159 ( .A(n91), .B(n92), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U160 ( .A(n87), .B(n88), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U161 ( .A(n81), .B(n82), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U162 ( .A(n79), .B(n80), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U163 ( .A(n77), .B(n78), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U164 ( .A(n62), .B(\b[0] ), .CI(n183), .CO(n61), .S(product[3]) );
  ADDFXL U165 ( .A(n121), .B(n122), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U166 ( .A(n71), .B(n72), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U167 ( .A(n83), .B(n84), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U168 ( .A(n75), .B(n76), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U169 ( .A(n65), .B(n66), .CI(n3), .CO(n2), .S(product[62]) );
  XNOR2XL U170 ( .A(b[61]), .B(b[60]), .Y(n322) );
  ADDFXL U171 ( .A(n69), .B(n70), .CI(n5), .CO(n4), .S(product[60]) );
  XOR2X1 U172 ( .A(n321), .B(n322), .Y(product[63]) );
  XOR2X1 U173 ( .A(n323), .B(b[63]), .Y(n321) );
  XNOR2X1 U174 ( .A(n64), .B(n2), .Y(n323) );
endmodule


module GSIM_DW01_add_499 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;
  assign SUM[0] = B[0];

  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2XL U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module GSIM_DW01_add_498 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module GSIM_DW01_add_497 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;

  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module GSIM_DW01_add_496 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;

  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  XOR3X2 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module GSIM_DW_mult_tc_3 ( a, b, product );
  input [3:0] a;
  input [63:0] b;
  output [67:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, \b[0] , \b[1] , n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318;
  assign product[1] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[2] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U3 ( .A(b[61]), .B(n317), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U4 ( .A(b[60]), .B(n316), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U5 ( .A(b[59]), .B(n315), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U6 ( .A(b[58]), .B(n314), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U7 ( .A(b[57]), .B(n313), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U8 ( .A(b[56]), .B(n312), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U9 ( .A(b[55]), .B(n311), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U10 ( .A(b[54]), .B(n310), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U11 ( .A(b[53]), .B(n309), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U12 ( .A(b[52]), .B(n308), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U13 ( .A(b[51]), .B(n307), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U14 ( .A(b[50]), .B(n306), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U15 ( .A(b[49]), .B(n305), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U16 ( .A(b[48]), .B(n304), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U17 ( .A(b[47]), .B(n303), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U18 ( .A(b[46]), .B(n302), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U19 ( .A(b[45]), .B(n301), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U20 ( .A(b[44]), .B(n300), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U21 ( .A(b[43]), .B(n299), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U22 ( .A(b[42]), .B(n298), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U23 ( .A(b[41]), .B(n297), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U24 ( .A(b[40]), .B(n296), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U25 ( .A(b[39]), .B(n295), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U26 ( .A(b[38]), .B(n294), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U27 ( .A(b[37]), .B(n293), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U28 ( .A(b[36]), .B(n292), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U29 ( .A(b[35]), .B(n291), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U30 ( .A(b[34]), .B(n290), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U31 ( .A(b[33]), .B(n289), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U32 ( .A(b[32]), .B(n288), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U33 ( .A(b[31]), .B(n287), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U34 ( .A(b[30]), .B(n286), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U35 ( .A(b[29]), .B(n285), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U36 ( .A(b[28]), .B(n284), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U37 ( .A(b[27]), .B(n283), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U38 ( .A(b[26]), .B(n282), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U39 ( .A(b[25]), .B(n281), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U40 ( .A(b[24]), .B(n280), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U41 ( .A(b[23]), .B(n279), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U42 ( .A(b[22]), .B(n278), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U43 ( .A(b[21]), .B(n277), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U44 ( .A(b[20]), .B(n276), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U45 ( .A(b[19]), .B(n275), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U46 ( .A(b[18]), .B(n274), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U47 ( .A(b[17]), .B(n273), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U48 ( .A(b[16]), .B(n272), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U49 ( .A(b[15]), .B(n271), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U50 ( .A(b[14]), .B(n270), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U51 ( .A(b[13]), .B(n269), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U52 ( .A(b[12]), .B(n268), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U53 ( .A(b[11]), .B(n267), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U54 ( .A(b[10]), .B(n266), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U55 ( .A(b[9]), .B(n265), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U56 ( .A(b[8]), .B(n264), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U57 ( .A(b[7]), .B(n263), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U58 ( .A(b[6]), .B(n262), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U59 ( .A(b[5]), .B(n261), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U60 ( .A(b[4]), .B(n260), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U61 ( .A(b[3]), .B(n259), .CI(n61), .CO(n60), .S(product[4]) );
  INVXL U131 ( .A(b[2]), .Y(n260) );
  XOR2XL U132 ( .A(b[2]), .B(\b[0] ), .Y(product[3]) );
  INVXL U133 ( .A(\b[1] ), .Y(n259) );
  XOR2XL U134 ( .A(n318), .B(b[60]), .Y(product[63]) );
  NAND2XL U135 ( .A(\b[0] ), .B(n260), .Y(n61) );
  INVXL U136 ( .A(b[12]), .Y(n270) );
  INVXL U137 ( .A(b[22]), .Y(n280) );
  INVXL U138 ( .A(b[32]), .Y(n290) );
  INVXL U139 ( .A(b[42]), .Y(n300) );
  INVXL U140 ( .A(b[52]), .Y(n310) );
  INVXL U141 ( .A(b[4]), .Y(n262) );
  INVXL U142 ( .A(b[3]), .Y(n261) );
  INVXL U143 ( .A(b[11]), .Y(n269) );
  INVXL U144 ( .A(b[21]), .Y(n279) );
  INVXL U145 ( .A(b[31]), .Y(n289) );
  INVXL U146 ( .A(b[41]), .Y(n299) );
  INVXL U147 ( .A(b[51]), .Y(n309) );
  INVXL U148 ( .A(b[14]), .Y(n272) );
  INVXL U149 ( .A(b[24]), .Y(n282) );
  INVXL U150 ( .A(b[34]), .Y(n292) );
  INVXL U151 ( .A(b[44]), .Y(n302) );
  INVXL U152 ( .A(b[54]), .Y(n312) );
  INVXL U153 ( .A(b[5]), .Y(n263) );
  INVXL U154 ( .A(b[6]), .Y(n264) );
  INVXL U155 ( .A(b[7]), .Y(n265) );
  INVXL U156 ( .A(b[8]), .Y(n266) );
  INVXL U157 ( .A(b[9]), .Y(n267) );
  INVXL U158 ( .A(b[10]), .Y(n268) );
  INVXL U159 ( .A(b[13]), .Y(n271) );
  INVXL U160 ( .A(b[15]), .Y(n273) );
  INVXL U161 ( .A(b[16]), .Y(n274) );
  INVXL U162 ( .A(b[17]), .Y(n275) );
  INVXL U163 ( .A(b[18]), .Y(n276) );
  INVXL U164 ( .A(b[19]), .Y(n277) );
  INVXL U165 ( .A(b[20]), .Y(n278) );
  INVXL U166 ( .A(b[23]), .Y(n281) );
  INVXL U167 ( .A(b[25]), .Y(n283) );
  INVXL U168 ( .A(b[26]), .Y(n284) );
  INVXL U169 ( .A(b[27]), .Y(n285) );
  INVXL U170 ( .A(b[28]), .Y(n286) );
  INVXL U171 ( .A(b[29]), .Y(n287) );
  INVXL U172 ( .A(b[30]), .Y(n288) );
  INVXL U173 ( .A(b[33]), .Y(n291) );
  INVXL U174 ( .A(b[35]), .Y(n293) );
  INVXL U175 ( .A(b[36]), .Y(n294) );
  INVXL U176 ( .A(b[37]), .Y(n295) );
  INVXL U177 ( .A(b[38]), .Y(n296) );
  INVXL U178 ( .A(b[39]), .Y(n297) );
  INVXL U179 ( .A(b[40]), .Y(n298) );
  INVXL U180 ( .A(b[43]), .Y(n301) );
  INVXL U181 ( .A(b[45]), .Y(n303) );
  INVXL U182 ( .A(b[46]), .Y(n304) );
  INVXL U183 ( .A(b[47]), .Y(n305) );
  INVXL U184 ( .A(b[48]), .Y(n306) );
  INVXL U185 ( .A(b[49]), .Y(n307) );
  INVXL U186 ( .A(b[50]), .Y(n308) );
  INVXL U187 ( .A(b[53]), .Y(n311) );
  INVXL U188 ( .A(b[55]), .Y(n313) );
  INVXL U189 ( .A(b[56]), .Y(n314) );
  INVXL U190 ( .A(b[57]), .Y(n315) );
  INVXL U191 ( .A(b[58]), .Y(n316) );
  INVXL U192 ( .A(b[59]), .Y(n317) );
  XNOR2X1 U193 ( .A(n2), .B(b[62]), .Y(n318) );
endmodule


module GSIM_DW_mult_tc_2 ( a, b, product );
  input [4:0] a;
  input [63:0] b;
  output [68:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, \b[0] , \b[1] , n321, n322, n323;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[1] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U4 ( .A(n67), .B(n68), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U6 ( .A(n71), .B(n72), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U12 ( .A(n83), .B(n84), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U14 ( .A(n87), .B(n88), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U16 ( .A(n91), .B(n92), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U18 ( .A(n95), .B(n96), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U20 ( .A(n99), .B(n100), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U22 ( .A(n103), .B(n104), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U24 ( .A(n107), .B(n108), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U26 ( .A(n111), .B(n112), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U28 ( .A(n115), .B(n116), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U30 ( .A(n119), .B(n120), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U50 ( .A(n159), .B(n160), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U52 ( .A(n163), .B(n164), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U54 ( .A(n167), .B(n168), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U56 ( .A(n171), .B(n172), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U58 ( .A(n175), .B(n176), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U60 ( .A(n179), .B(n180), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U62 ( .A(n62), .B(\b[0] ), .CI(n183), .CO(n61), .S(product[3]) );
  ADDHXL U63 ( .A(\b[0] ), .B(b[2]), .CO(n62), .S(product[2]) );
  ADDFXL U65 ( .A(b[59]), .B(b[62]), .CI(b[60]), .CO(n64), .S(n65) );
  ADDFXL U66 ( .A(b[58]), .B(b[61]), .CI(b[59]), .CO(n66), .S(n67) );
  ADDFXL U67 ( .A(b[57]), .B(b[60]), .CI(b[58]), .CO(n68), .S(n69) );
  ADDFXL U68 ( .A(b[56]), .B(b[59]), .CI(b[57]), .CO(n70), .S(n71) );
  ADDFXL U69 ( .A(b[55]), .B(b[58]), .CI(b[56]), .CO(n72), .S(n73) );
  ADDFXL U70 ( .A(b[54]), .B(b[57]), .CI(b[55]), .CO(n74), .S(n75) );
  ADDFXL U71 ( .A(b[53]), .B(b[56]), .CI(b[54]), .CO(n76), .S(n77) );
  ADDFXL U72 ( .A(b[52]), .B(b[55]), .CI(b[53]), .CO(n78), .S(n79) );
  ADDFXL U73 ( .A(b[51]), .B(b[54]), .CI(b[52]), .CO(n80), .S(n81) );
  ADDFXL U74 ( .A(b[50]), .B(b[53]), .CI(b[51]), .CO(n82), .S(n83) );
  ADDFXL U75 ( .A(b[49]), .B(b[52]), .CI(b[50]), .CO(n84), .S(n85) );
  ADDFXL U76 ( .A(b[48]), .B(b[51]), .CI(b[49]), .CO(n86), .S(n87) );
  ADDFXL U77 ( .A(b[47]), .B(b[50]), .CI(b[48]), .CO(n88), .S(n89) );
  ADDFXL U78 ( .A(b[46]), .B(b[49]), .CI(b[47]), .CO(n90), .S(n91) );
  ADDFXL U79 ( .A(b[45]), .B(b[48]), .CI(b[46]), .CO(n92), .S(n93) );
  ADDFXL U80 ( .A(b[44]), .B(b[47]), .CI(b[45]), .CO(n94), .S(n95) );
  ADDFXL U81 ( .A(b[43]), .B(b[46]), .CI(b[44]), .CO(n96), .S(n97) );
  ADDFXL U82 ( .A(b[42]), .B(b[45]), .CI(b[43]), .CO(n98), .S(n99) );
  ADDFXL U83 ( .A(b[41]), .B(b[44]), .CI(b[42]), .CO(n100), .S(n101) );
  ADDFXL U84 ( .A(b[40]), .B(b[43]), .CI(b[41]), .CO(n102), .S(n103) );
  ADDFXL U85 ( .A(b[39]), .B(b[42]), .CI(b[40]), .CO(n104), .S(n105) );
  ADDFXL U86 ( .A(b[38]), .B(b[41]), .CI(b[39]), .CO(n106), .S(n107) );
  ADDFXL U87 ( .A(b[37]), .B(b[40]), .CI(b[38]), .CO(n108), .S(n109) );
  ADDFXL U88 ( .A(b[36]), .B(b[39]), .CI(b[37]), .CO(n110), .S(n111) );
  ADDFXL U89 ( .A(b[35]), .B(b[38]), .CI(b[36]), .CO(n112), .S(n113) );
  ADDFXL U90 ( .A(b[34]), .B(b[37]), .CI(b[35]), .CO(n114), .S(n115) );
  ADDFXL U91 ( .A(b[33]), .B(b[36]), .CI(b[34]), .CO(n116), .S(n117) );
  ADDFXL U92 ( .A(b[32]), .B(b[35]), .CI(b[33]), .CO(n118), .S(n119) );
  ADDFXL U93 ( .A(b[31]), .B(b[34]), .CI(b[32]), .CO(n120), .S(n121) );
  ADDFXL U94 ( .A(b[30]), .B(b[33]), .CI(b[31]), .CO(n122), .S(n123) );
  ADDFXL U95 ( .A(b[29]), .B(b[32]), .CI(b[30]), .CO(n124), .S(n125) );
  ADDFXL U96 ( .A(b[28]), .B(b[31]), .CI(b[29]), .CO(n126), .S(n127) );
  ADDFXL U97 ( .A(b[27]), .B(b[30]), .CI(b[28]), .CO(n128), .S(n129) );
  ADDFXL U98 ( .A(b[26]), .B(b[29]), .CI(b[27]), .CO(n130), .S(n131) );
  ADDFXL U99 ( .A(b[25]), .B(b[28]), .CI(b[26]), .CO(n132), .S(n133) );
  ADDFXL U100 ( .A(b[24]), .B(b[27]), .CI(b[25]), .CO(n134), .S(n135) );
  ADDFXL U101 ( .A(b[23]), .B(b[26]), .CI(b[24]), .CO(n136), .S(n137) );
  ADDFXL U102 ( .A(b[22]), .B(b[25]), .CI(b[23]), .CO(n138), .S(n139) );
  ADDFXL U103 ( .A(b[21]), .B(b[24]), .CI(b[22]), .CO(n140), .S(n141) );
  ADDFXL U104 ( .A(b[20]), .B(b[23]), .CI(b[21]), .CO(n142), .S(n143) );
  ADDFXL U105 ( .A(b[19]), .B(b[22]), .CI(b[20]), .CO(n144), .S(n145) );
  ADDFXL U106 ( .A(b[18]), .B(b[21]), .CI(b[19]), .CO(n146), .S(n147) );
  ADDFXL U107 ( .A(b[17]), .B(b[20]), .CI(b[18]), .CO(n148), .S(n149) );
  ADDFXL U108 ( .A(b[16]), .B(b[19]), .CI(b[17]), .CO(n150), .S(n151) );
  ADDFXL U109 ( .A(b[15]), .B(b[18]), .CI(b[16]), .CO(n152), .S(n153) );
  ADDFXL U110 ( .A(b[14]), .B(b[17]), .CI(b[15]), .CO(n154), .S(n155) );
  ADDFXL U111 ( .A(b[13]), .B(b[16]), .CI(b[14]), .CO(n156), .S(n157) );
  ADDFXL U112 ( .A(b[12]), .B(b[15]), .CI(b[13]), .CO(n158), .S(n159) );
  ADDFXL U113 ( .A(b[11]), .B(b[14]), .CI(b[12]), .CO(n160), .S(n161) );
  ADDFXL U114 ( .A(b[10]), .B(b[13]), .CI(b[11]), .CO(n162), .S(n163) );
  ADDFXL U115 ( .A(b[9]), .B(b[12]), .CI(b[10]), .CO(n164), .S(n165) );
  ADDFXL U116 ( .A(b[8]), .B(b[11]), .CI(b[9]), .CO(n166), .S(n167) );
  ADDFXL U117 ( .A(b[7]), .B(b[10]), .CI(b[8]), .CO(n168), .S(n169) );
  ADDFXL U118 ( .A(b[6]), .B(b[9]), .CI(b[7]), .CO(n170), .S(n171) );
  ADDFXL U119 ( .A(b[5]), .B(b[8]), .CI(b[6]), .CO(n172), .S(n173) );
  ADDFXL U121 ( .A(b[3]), .B(b[6]), .CI(b[4]), .CO(n176), .S(n177) );
  ADDFXL U122 ( .A(b[2]), .B(b[5]), .CI(b[3]), .CO(n178), .S(n179) );
  ADDHXL U124 ( .A(b[3]), .B(\b[1] ), .CO(n182), .S(n183) );
  ADDFXL U129 ( .A(n161), .B(n162), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U130 ( .A(n157), .B(n158), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U131 ( .A(n155), .B(n156), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U132 ( .A(n153), .B(n154), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U133 ( .A(n151), .B(n152), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U134 ( .A(n149), .B(n150), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U135 ( .A(n147), .B(n148), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U136 ( .A(n139), .B(n140), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U137 ( .A(n141), .B(n142), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U138 ( .A(n143), .B(n144), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U139 ( .A(n145), .B(n146), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U140 ( .A(\b[1] ), .B(b[4]), .CI(b[2]), .CO(n180), .S(n181) );
  ADDFXL U141 ( .A(n165), .B(n166), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U142 ( .A(n169), .B(n170), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U143 ( .A(n137), .B(n138), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U144 ( .A(n135), .B(n136), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U145 ( .A(n133), .B(n134), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U146 ( .A(n131), .B(n132), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U147 ( .A(n129), .B(n130), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U148 ( .A(n127), .B(n128), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U149 ( .A(n125), .B(n126), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U150 ( .A(n121), .B(n122), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U151 ( .A(n117), .B(n118), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U152 ( .A(n113), .B(n114), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U153 ( .A(n109), .B(n110), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U154 ( .A(n105), .B(n106), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U155 ( .A(n101), .B(n102), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U156 ( .A(n97), .B(n98), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U157 ( .A(n93), .B(n94), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U158 ( .A(n89), .B(n90), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U159 ( .A(n85), .B(n86), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U160 ( .A(n81), .B(n82), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U161 ( .A(n79), .B(n80), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U162 ( .A(n77), .B(n78), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U163 ( .A(n75), .B(n76), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U164 ( .A(n73), .B(n74), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U165 ( .A(n123), .B(n124), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U166 ( .A(n181), .B(n182), .CI(n61), .CO(n60), .S(product[4]) );
  ADDFXL U167 ( .A(n69), .B(n70), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U168 ( .A(n177), .B(n178), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U169 ( .A(n173), .B(n174), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U170 ( .A(n65), .B(n66), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U171 ( .A(b[4]), .B(b[7]), .CI(b[5]), .CO(n174), .S(n175) );
  XNOR2XL U172 ( .A(b[61]), .B(b[60]), .Y(n322) );
  XOR2X1 U173 ( .A(n321), .B(n322), .Y(product[63]) );
  XOR2X1 U174 ( .A(n323), .B(b[63]), .Y(n321) );
  XNOR2X1 U175 ( .A(n64), .B(n2), .Y(n323) );
endmodule


module GSIM_DW_mult_tc_1 ( a, b, product );
  input [4:0] a;
  input [63:0] b;
  output [68:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, \b[0] , \b[1] , n321, n322, n323;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[1] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U4 ( .A(n67), .B(n68), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U5 ( .A(n69), .B(n70), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U14 ( .A(n87), .B(n88), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U16 ( .A(n91), .B(n92), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U20 ( .A(n99), .B(n100), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U22 ( .A(n103), .B(n104), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U24 ( .A(n107), .B(n108), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U26 ( .A(n111), .B(n112), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U28 ( .A(n115), .B(n116), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U30 ( .A(n119), .B(n120), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U52 ( .A(n163), .B(n164), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U54 ( .A(n167), .B(n168), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U56 ( .A(n171), .B(n172), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U58 ( .A(n175), .B(n176), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U60 ( .A(n179), .B(n180), .CI(n60), .CO(n59), .S(product[5]) );
  ADDHXL U63 ( .A(\b[0] ), .B(b[2]), .CO(n62), .S(product[2]) );
  ADDFXL U65 ( .A(b[59]), .B(b[62]), .CI(b[60]), .CO(n64), .S(n65) );
  ADDFXL U66 ( .A(b[58]), .B(b[61]), .CI(b[59]), .CO(n66), .S(n67) );
  ADDFXL U67 ( .A(b[57]), .B(b[60]), .CI(b[58]), .CO(n68), .S(n69) );
  ADDFXL U68 ( .A(b[56]), .B(b[59]), .CI(b[57]), .CO(n70), .S(n71) );
  ADDFXL U69 ( .A(b[55]), .B(b[58]), .CI(b[56]), .CO(n72), .S(n73) );
  ADDFXL U70 ( .A(b[54]), .B(b[57]), .CI(b[55]), .CO(n74), .S(n75) );
  ADDFXL U71 ( .A(b[53]), .B(b[56]), .CI(b[54]), .CO(n76), .S(n77) );
  ADDFXL U72 ( .A(b[52]), .B(b[55]), .CI(b[53]), .CO(n78), .S(n79) );
  ADDFXL U73 ( .A(b[51]), .B(b[54]), .CI(b[52]), .CO(n80), .S(n81) );
  ADDFXL U74 ( .A(b[50]), .B(b[53]), .CI(b[51]), .CO(n82), .S(n83) );
  ADDFXL U75 ( .A(b[49]), .B(b[52]), .CI(b[50]), .CO(n84), .S(n85) );
  ADDFXL U76 ( .A(b[48]), .B(b[51]), .CI(b[49]), .CO(n86), .S(n87) );
  ADDFXL U77 ( .A(b[47]), .B(b[50]), .CI(b[48]), .CO(n88), .S(n89) );
  ADDFXL U78 ( .A(b[46]), .B(b[49]), .CI(b[47]), .CO(n90), .S(n91) );
  ADDFXL U79 ( .A(b[45]), .B(b[48]), .CI(b[46]), .CO(n92), .S(n93) );
  ADDFXL U80 ( .A(b[44]), .B(b[47]), .CI(b[45]), .CO(n94), .S(n95) );
  ADDFXL U81 ( .A(b[43]), .B(b[46]), .CI(b[44]), .CO(n96), .S(n97) );
  ADDFXL U82 ( .A(b[42]), .B(b[45]), .CI(b[43]), .CO(n98), .S(n99) );
  ADDFXL U83 ( .A(b[41]), .B(b[44]), .CI(b[42]), .CO(n100), .S(n101) );
  ADDFXL U84 ( .A(b[40]), .B(b[43]), .CI(b[41]), .CO(n102), .S(n103) );
  ADDFXL U85 ( .A(b[39]), .B(b[42]), .CI(b[40]), .CO(n104), .S(n105) );
  ADDFXL U86 ( .A(b[38]), .B(b[41]), .CI(b[39]), .CO(n106), .S(n107) );
  ADDFXL U87 ( .A(b[37]), .B(b[40]), .CI(b[38]), .CO(n108), .S(n109) );
  ADDFXL U88 ( .A(b[36]), .B(b[39]), .CI(b[37]), .CO(n110), .S(n111) );
  ADDFXL U89 ( .A(b[35]), .B(b[38]), .CI(b[36]), .CO(n112), .S(n113) );
  ADDFXL U90 ( .A(b[34]), .B(b[37]), .CI(b[35]), .CO(n114), .S(n115) );
  ADDFXL U91 ( .A(b[33]), .B(b[36]), .CI(b[34]), .CO(n116), .S(n117) );
  ADDFXL U92 ( .A(b[32]), .B(b[35]), .CI(b[33]), .CO(n118), .S(n119) );
  ADDFXL U93 ( .A(b[31]), .B(b[34]), .CI(b[32]), .CO(n120), .S(n121) );
  ADDFXL U94 ( .A(b[30]), .B(b[33]), .CI(b[31]), .CO(n122), .S(n123) );
  ADDFXL U95 ( .A(b[29]), .B(b[32]), .CI(b[30]), .CO(n124), .S(n125) );
  ADDFXL U96 ( .A(b[28]), .B(b[31]), .CI(b[29]), .CO(n126), .S(n127) );
  ADDFXL U97 ( .A(b[27]), .B(b[30]), .CI(b[28]), .CO(n128), .S(n129) );
  ADDFXL U98 ( .A(b[26]), .B(b[29]), .CI(b[27]), .CO(n130), .S(n131) );
  ADDFXL U99 ( .A(b[25]), .B(b[28]), .CI(b[26]), .CO(n132), .S(n133) );
  ADDFXL U100 ( .A(b[24]), .B(b[27]), .CI(b[25]), .CO(n134), .S(n135) );
  ADDFXL U101 ( .A(b[23]), .B(b[26]), .CI(b[24]), .CO(n136), .S(n137) );
  ADDFXL U102 ( .A(b[22]), .B(b[25]), .CI(b[23]), .CO(n138), .S(n139) );
  ADDFXL U103 ( .A(b[21]), .B(b[24]), .CI(b[22]), .CO(n140), .S(n141) );
  ADDFXL U104 ( .A(b[20]), .B(b[23]), .CI(b[21]), .CO(n142), .S(n143) );
  ADDFXL U105 ( .A(b[19]), .B(b[22]), .CI(b[20]), .CO(n144), .S(n145) );
  ADDFXL U106 ( .A(b[18]), .B(b[21]), .CI(b[19]), .CO(n146), .S(n147) );
  ADDFXL U107 ( .A(b[17]), .B(b[20]), .CI(b[18]), .CO(n148), .S(n149) );
  ADDFXL U108 ( .A(b[16]), .B(b[19]), .CI(b[17]), .CO(n150), .S(n151) );
  ADDFXL U109 ( .A(b[15]), .B(b[18]), .CI(b[16]), .CO(n152), .S(n153) );
  ADDFXL U110 ( .A(b[14]), .B(b[17]), .CI(b[15]), .CO(n154), .S(n155) );
  ADDFXL U111 ( .A(b[13]), .B(b[16]), .CI(b[14]), .CO(n156), .S(n157) );
  ADDFXL U112 ( .A(b[12]), .B(b[15]), .CI(b[13]), .CO(n158), .S(n159) );
  ADDFXL U113 ( .A(b[11]), .B(b[14]), .CI(b[12]), .CO(n160), .S(n161) );
  ADDFXL U114 ( .A(b[10]), .B(b[13]), .CI(b[11]), .CO(n162), .S(n163) );
  ADDFXL U115 ( .A(b[9]), .B(b[12]), .CI(b[10]), .CO(n164), .S(n165) );
  ADDFXL U116 ( .A(b[8]), .B(b[11]), .CI(b[9]), .CO(n166), .S(n167) );
  ADDFXL U117 ( .A(b[7]), .B(b[10]), .CI(b[8]), .CO(n168), .S(n169) );
  ADDFXL U118 ( .A(b[6]), .B(b[9]), .CI(b[7]), .CO(n170), .S(n171) );
  ADDFXL U119 ( .A(b[5]), .B(b[8]), .CI(b[6]), .CO(n172), .S(n173) );
  ADDFXL U120 ( .A(b[4]), .B(b[7]), .CI(b[5]), .CO(n174), .S(n175) );
  ADDFXL U121 ( .A(b[3]), .B(b[6]), .CI(b[4]), .CO(n176), .S(n177) );
  ADDFXL U123 ( .A(\b[1] ), .B(b[4]), .CI(b[2]), .CO(n180), .S(n181) );
  ADDHXL U124 ( .A(b[3]), .B(\b[1] ), .CO(n182), .S(n183) );
  ADDFXL U129 ( .A(b[2]), .B(b[5]), .CI(b[3]), .CO(n178), .S(n179) );
  ADDFXL U130 ( .A(n161), .B(n162), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U131 ( .A(n157), .B(n158), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U132 ( .A(n159), .B(n160), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U133 ( .A(n155), .B(n156), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U134 ( .A(n153), .B(n154), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U135 ( .A(n151), .B(n152), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U136 ( .A(n149), .B(n150), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U137 ( .A(n147), .B(n148), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U138 ( .A(n139), .B(n140), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U139 ( .A(n141), .B(n142), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U140 ( .A(n143), .B(n144), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U141 ( .A(n145), .B(n146), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U142 ( .A(n165), .B(n166), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U143 ( .A(n169), .B(n170), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U144 ( .A(n173), .B(n174), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U145 ( .A(n177), .B(n178), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U146 ( .A(n137), .B(n138), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U147 ( .A(n135), .B(n136), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U148 ( .A(n133), .B(n134), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U149 ( .A(n131), .B(n132), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U150 ( .A(n129), .B(n130), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U151 ( .A(n127), .B(n128), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U152 ( .A(n125), .B(n126), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U153 ( .A(n121), .B(n122), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U154 ( .A(n117), .B(n118), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U155 ( .A(n113), .B(n114), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U156 ( .A(n109), .B(n110), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U157 ( .A(n105), .B(n106), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U158 ( .A(n101), .B(n102), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U159 ( .A(n97), .B(n98), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U160 ( .A(n93), .B(n94), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U161 ( .A(n89), .B(n90), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U162 ( .A(n85), .B(n86), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U163 ( .A(n83), .B(n84), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U164 ( .A(n81), .B(n82), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U165 ( .A(n79), .B(n80), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U166 ( .A(n77), .B(n78), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U167 ( .A(n75), .B(n76), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U168 ( .A(n181), .B(n182), .CI(n61), .CO(n60), .S(product[4]) );
  ADDFXL U169 ( .A(n62), .B(\b[0] ), .CI(n183), .CO(n61), .S(product[3]) );
  ADDFXL U170 ( .A(n71), .B(n72), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U171 ( .A(n65), .B(n66), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U172 ( .A(n123), .B(n124), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U173 ( .A(n73), .B(n74), .CI(n7), .CO(n6), .S(product[58]) );
  XNOR2XL U174 ( .A(b[61]), .B(b[60]), .Y(n322) );
  ADDFXL U175 ( .A(n95), .B(n96), .CI(n18), .CO(n17), .S(product[47]) );
  XOR2X1 U176 ( .A(n321), .B(n322), .Y(product[63]) );
  XOR2X1 U177 ( .A(n323), .B(b[63]), .Y(n321) );
  XNOR2X1 U178 ( .A(n64), .B(n2), .Y(n323) );
endmodule


module GSIM_DW_mult_tc_0 ( a, b, product );
  input [3:0] a;
  input [63:0] b;
  output [67:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, \b[0] , \b[1] , n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318;
  assign product[1] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[2] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U3 ( .A(b[61]), .B(n317), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U4 ( .A(b[60]), .B(n316), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U5 ( .A(b[59]), .B(n315), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U6 ( .A(b[58]), .B(n314), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U7 ( .A(b[57]), .B(n313), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U8 ( .A(b[56]), .B(n312), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U9 ( .A(b[55]), .B(n311), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U10 ( .A(b[54]), .B(n310), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U11 ( .A(b[53]), .B(n309), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U12 ( .A(b[52]), .B(n308), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U13 ( .A(b[51]), .B(n307), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U14 ( .A(b[50]), .B(n306), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U15 ( .A(b[49]), .B(n305), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U16 ( .A(b[48]), .B(n304), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U17 ( .A(b[47]), .B(n303), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U18 ( .A(b[46]), .B(n302), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U19 ( .A(b[45]), .B(n301), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U20 ( .A(b[44]), .B(n300), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U21 ( .A(b[43]), .B(n299), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U22 ( .A(b[42]), .B(n298), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U23 ( .A(b[41]), .B(n297), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U24 ( .A(b[40]), .B(n296), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U25 ( .A(b[39]), .B(n295), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U26 ( .A(b[38]), .B(n294), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U27 ( .A(b[37]), .B(n293), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U28 ( .A(b[36]), .B(n292), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U29 ( .A(b[35]), .B(n291), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U30 ( .A(b[34]), .B(n290), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U31 ( .A(b[33]), .B(n289), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U32 ( .A(b[32]), .B(n288), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U33 ( .A(b[31]), .B(n287), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U34 ( .A(b[30]), .B(n286), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U35 ( .A(b[29]), .B(n285), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U36 ( .A(b[28]), .B(n284), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U37 ( .A(b[27]), .B(n283), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U38 ( .A(b[26]), .B(n282), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U39 ( .A(b[25]), .B(n281), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U40 ( .A(b[24]), .B(n280), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U41 ( .A(b[23]), .B(n279), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U42 ( .A(b[22]), .B(n278), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U43 ( .A(b[21]), .B(n277), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U44 ( .A(b[20]), .B(n276), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U45 ( .A(b[19]), .B(n275), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U46 ( .A(b[18]), .B(n274), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U47 ( .A(b[17]), .B(n273), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U48 ( .A(b[16]), .B(n272), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U49 ( .A(b[15]), .B(n271), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U50 ( .A(b[14]), .B(n270), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U51 ( .A(b[13]), .B(n269), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U52 ( .A(b[12]), .B(n268), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U53 ( .A(b[11]), .B(n267), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U54 ( .A(b[10]), .B(n266), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U55 ( .A(b[9]), .B(n265), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U56 ( .A(b[8]), .B(n264), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U57 ( .A(b[7]), .B(n263), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U58 ( .A(b[6]), .B(n262), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U59 ( .A(b[5]), .B(n261), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U60 ( .A(b[4]), .B(n260), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U61 ( .A(b[3]), .B(n259), .CI(n61), .CO(n60), .S(product[4]) );
  NAND2XL U131 ( .A(\b[0] ), .B(n260), .Y(n61) );
  INVXL U132 ( .A(\b[1] ), .Y(n259) );
  INVXL U133 ( .A(b[18]), .Y(n276) );
  INVXL U134 ( .A(b[28]), .Y(n286) );
  INVXL U135 ( .A(b[38]), .Y(n296) );
  INVXL U136 ( .A(b[48]), .Y(n306) );
  INVXL U137 ( .A(b[10]), .Y(n268) );
  INVXL U138 ( .A(b[17]), .Y(n275) );
  INVXL U139 ( .A(b[19]), .Y(n277) );
  INVXL U140 ( .A(b[20]), .Y(n278) );
  INVXL U141 ( .A(b[27]), .Y(n285) );
  INVXL U142 ( .A(b[29]), .Y(n287) );
  INVXL U143 ( .A(b[30]), .Y(n288) );
  INVXL U144 ( .A(b[37]), .Y(n295) );
  INVXL U145 ( .A(b[39]), .Y(n297) );
  INVXL U146 ( .A(b[40]), .Y(n298) );
  INVXL U147 ( .A(b[47]), .Y(n305) );
  INVXL U148 ( .A(b[49]), .Y(n307) );
  INVXL U149 ( .A(b[50]), .Y(n308) );
  INVXL U150 ( .A(b[51]), .Y(n309) );
  INVXL U151 ( .A(b[6]), .Y(n264) );
  INVXL U152 ( .A(b[7]), .Y(n265) );
  INVXL U153 ( .A(b[8]), .Y(n266) );
  INVXL U154 ( .A(b[9]), .Y(n267) );
  INVXL U155 ( .A(b[16]), .Y(n274) );
  INVXL U156 ( .A(b[26]), .Y(n284) );
  INVXL U157 ( .A(b[36]), .Y(n294) );
  INVXL U158 ( .A(b[46]), .Y(n304) );
  INVXL U159 ( .A(b[3]), .Y(n261) );
  INVXL U160 ( .A(b[4]), .Y(n262) );
  INVXL U161 ( .A(b[5]), .Y(n263) );
  INVXL U162 ( .A(b[11]), .Y(n269) );
  INVXL U163 ( .A(b[12]), .Y(n270) );
  INVXL U164 ( .A(b[13]), .Y(n271) );
  INVXL U165 ( .A(b[14]), .Y(n272) );
  INVXL U166 ( .A(b[15]), .Y(n273) );
  INVXL U167 ( .A(b[21]), .Y(n279) );
  INVXL U168 ( .A(b[22]), .Y(n280) );
  INVXL U169 ( .A(b[23]), .Y(n281) );
  INVXL U170 ( .A(b[24]), .Y(n282) );
  INVXL U171 ( .A(b[25]), .Y(n283) );
  INVXL U172 ( .A(b[31]), .Y(n289) );
  INVXL U173 ( .A(b[32]), .Y(n290) );
  INVXL U174 ( .A(b[33]), .Y(n291) );
  INVXL U175 ( .A(b[34]), .Y(n292) );
  INVXL U176 ( .A(b[35]), .Y(n293) );
  INVXL U177 ( .A(b[41]), .Y(n299) );
  INVXL U178 ( .A(b[42]), .Y(n300) );
  INVXL U179 ( .A(b[43]), .Y(n301) );
  INVXL U180 ( .A(b[44]), .Y(n302) );
  INVXL U181 ( .A(b[45]), .Y(n303) );
  INVXL U182 ( .A(b[52]), .Y(n310) );
  INVXL U183 ( .A(b[53]), .Y(n311) );
  INVXL U184 ( .A(b[54]), .Y(n312) );
  INVXL U185 ( .A(b[55]), .Y(n313) );
  INVXL U186 ( .A(b[56]), .Y(n314) );
  INVXL U187 ( .A(b[57]), .Y(n315) );
  INVXL U188 ( .A(b[58]), .Y(n316) );
  INVXL U189 ( .A(b[59]), .Y(n317) );
  INVXL U190 ( .A(b[2]), .Y(n260) );
  XOR2X1 U191 ( .A(n318), .B(b[60]), .Y(product[63]) );
  XNOR2X1 U192 ( .A(n2), .B(b[62]), .Y(n318) );
  XOR2X1 U193 ( .A(b[2]), .B(\b[0] ), .Y(product[3]) );
endmodule


module GSIM_DW01_add_476 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;
  assign SUM[0] = B[0];

  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module GSIM_DW01_add_475 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;
  assign SUM[15] = B[15];
  assign SUM[14] = B[14];
  assign SUM[13] = B[13];
  assign SUM[12] = B[12];
  assign SUM[11] = B[11];
  assign SUM[10] = B[10];
  assign SUM[9] = B[9];
  assign SUM[8] = B[8];
  assign SUM[7] = B[7];
  assign SUM[6] = B[6];
  assign SUM[5] = B[5];
  assign SUM[4] = B[4];
  assign SUM[3] = B[3];
  assign SUM[2] = B[2];
  assign SUM[1] = B[1];

  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(n1), .CO(carry[18]), .S(SUM[17]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  AND2X2 U1 ( .A(B[16]), .B(A[16]), .Y(n1) );
  XOR2XL U2 ( .A(B[16]), .B(A[16]), .Y(SUM[16]) );
endmodule


module GSIM_DW01_add_474 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;
  assign SUM[0] = A[0];

  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2XL U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module GSIM_DW01_add_473 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module GSIM_DW01_add_472 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  XOR3X2 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module GSIM_DW_mult_tc_8 ( a, b, product );
  input [4:0] a;
  input [63:0] b;
  output [68:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, \b[0] , \b[1] , n321, n322, n323;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[1] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U4 ( .A(n67), .B(n68), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U5 ( .A(n69), .B(n70), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U12 ( .A(n83), .B(n84), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U16 ( .A(n91), .B(n92), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U18 ( .A(n95), .B(n96), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U20 ( .A(n99), .B(n100), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U46 ( .A(n151), .B(n152), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U48 ( .A(n155), .B(n156), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U50 ( .A(n159), .B(n160), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U52 ( .A(n163), .B(n164), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U56 ( .A(n171), .B(n172), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U58 ( .A(n175), .B(n176), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U60 ( .A(n179), .B(n180), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U65 ( .A(b[59]), .B(b[62]), .CI(b[60]), .CO(n64), .S(n65) );
  ADDFXL U66 ( .A(b[58]), .B(b[61]), .CI(b[59]), .CO(n66), .S(n67) );
  ADDFXL U67 ( .A(b[57]), .B(b[60]), .CI(b[58]), .CO(n68), .S(n69) );
  ADDFXL U68 ( .A(b[56]), .B(b[59]), .CI(b[57]), .CO(n70), .S(n71) );
  ADDFXL U69 ( .A(b[55]), .B(b[58]), .CI(b[56]), .CO(n72), .S(n73) );
  ADDFXL U70 ( .A(b[54]), .B(b[57]), .CI(b[55]), .CO(n74), .S(n75) );
  ADDFXL U71 ( .A(b[53]), .B(b[56]), .CI(b[54]), .CO(n76), .S(n77) );
  ADDFXL U72 ( .A(b[52]), .B(b[55]), .CI(b[53]), .CO(n78), .S(n79) );
  ADDFXL U73 ( .A(b[51]), .B(b[54]), .CI(b[52]), .CO(n80), .S(n81) );
  ADDFXL U74 ( .A(b[50]), .B(b[53]), .CI(b[51]), .CO(n82), .S(n83) );
  ADDFXL U75 ( .A(b[49]), .B(b[52]), .CI(b[50]), .CO(n84), .S(n85) );
  ADDFXL U76 ( .A(b[48]), .B(b[51]), .CI(b[49]), .CO(n86), .S(n87) );
  ADDFXL U77 ( .A(b[47]), .B(b[50]), .CI(b[48]), .CO(n88), .S(n89) );
  ADDFXL U78 ( .A(b[46]), .B(b[49]), .CI(b[47]), .CO(n90), .S(n91) );
  ADDFXL U79 ( .A(b[45]), .B(b[48]), .CI(b[46]), .CO(n92), .S(n93) );
  ADDFXL U80 ( .A(b[44]), .B(b[47]), .CI(b[45]), .CO(n94), .S(n95) );
  ADDFXL U81 ( .A(b[43]), .B(b[46]), .CI(b[44]), .CO(n96), .S(n97) );
  ADDFXL U82 ( .A(b[42]), .B(b[45]), .CI(b[43]), .CO(n98), .S(n99) );
  ADDFXL U83 ( .A(b[41]), .B(b[44]), .CI(b[42]), .CO(n100), .S(n101) );
  ADDFXL U84 ( .A(b[40]), .B(b[43]), .CI(b[41]), .CO(n102), .S(n103) );
  ADDFXL U85 ( .A(b[39]), .B(b[42]), .CI(b[40]), .CO(n104), .S(n105) );
  ADDFXL U86 ( .A(b[38]), .B(b[41]), .CI(b[39]), .CO(n106), .S(n107) );
  ADDFXL U87 ( .A(b[37]), .B(b[40]), .CI(b[38]), .CO(n108), .S(n109) );
  ADDFXL U88 ( .A(b[36]), .B(b[39]), .CI(b[37]), .CO(n110), .S(n111) );
  ADDFXL U89 ( .A(b[35]), .B(b[38]), .CI(b[36]), .CO(n112), .S(n113) );
  ADDFXL U90 ( .A(b[34]), .B(b[37]), .CI(b[35]), .CO(n114), .S(n115) );
  ADDFXL U91 ( .A(b[33]), .B(b[36]), .CI(b[34]), .CO(n116), .S(n117) );
  ADDFXL U92 ( .A(b[32]), .B(b[35]), .CI(b[33]), .CO(n118), .S(n119) );
  ADDFXL U93 ( .A(b[31]), .B(b[34]), .CI(b[32]), .CO(n120), .S(n121) );
  ADDFXL U94 ( .A(b[30]), .B(b[33]), .CI(b[31]), .CO(n122), .S(n123) );
  ADDFXL U95 ( .A(b[29]), .B(b[32]), .CI(b[30]), .CO(n124), .S(n125) );
  ADDFXL U96 ( .A(b[28]), .B(b[31]), .CI(b[29]), .CO(n126), .S(n127) );
  ADDFXL U97 ( .A(b[27]), .B(b[30]), .CI(b[28]), .CO(n128), .S(n129) );
  ADDFXL U98 ( .A(b[26]), .B(b[29]), .CI(b[27]), .CO(n130), .S(n131) );
  ADDFXL U99 ( .A(b[25]), .B(b[28]), .CI(b[26]), .CO(n132), .S(n133) );
  ADDFXL U100 ( .A(b[24]), .B(b[27]), .CI(b[25]), .CO(n134), .S(n135) );
  ADDFXL U101 ( .A(b[23]), .B(b[26]), .CI(b[24]), .CO(n136), .S(n137) );
  ADDFXL U102 ( .A(b[22]), .B(b[25]), .CI(b[23]), .CO(n138), .S(n139) );
  ADDFXL U103 ( .A(b[21]), .B(b[24]), .CI(b[22]), .CO(n140), .S(n141) );
  ADDFXL U104 ( .A(b[20]), .B(b[23]), .CI(b[21]), .CO(n142), .S(n143) );
  ADDFXL U105 ( .A(b[19]), .B(b[22]), .CI(b[20]), .CO(n144), .S(n145) );
  ADDFXL U106 ( .A(b[18]), .B(b[21]), .CI(b[19]), .CO(n146), .S(n147) );
  ADDFXL U107 ( .A(b[17]), .B(b[20]), .CI(b[18]), .CO(n148), .S(n149) );
  ADDFXL U108 ( .A(b[16]), .B(b[19]), .CI(b[17]), .CO(n150), .S(n151) );
  ADDFXL U109 ( .A(b[15]), .B(b[18]), .CI(b[16]), .CO(n152), .S(n153) );
  ADDFXL U110 ( .A(b[14]), .B(b[17]), .CI(b[15]), .CO(n154), .S(n155) );
  ADDFXL U111 ( .A(b[13]), .B(b[16]), .CI(b[14]), .CO(n156), .S(n157) );
  ADDFXL U112 ( .A(b[12]), .B(b[15]), .CI(b[13]), .CO(n158), .S(n159) );
  ADDFXL U113 ( .A(b[11]), .B(b[14]), .CI(b[12]), .CO(n160), .S(n161) );
  ADDFXL U114 ( .A(b[10]), .B(b[13]), .CI(b[11]), .CO(n162), .S(n163) );
  ADDFXL U115 ( .A(b[9]), .B(b[12]), .CI(b[10]), .CO(n164), .S(n165) );
  ADDFXL U116 ( .A(b[8]), .B(b[11]), .CI(b[9]), .CO(n166), .S(n167) );
  ADDFXL U117 ( .A(b[7]), .B(b[10]), .CI(b[8]), .CO(n168), .S(n169) );
  ADDFXL U118 ( .A(b[6]), .B(b[9]), .CI(b[7]), .CO(n170), .S(n171) );
  ADDFXL U119 ( .A(b[5]), .B(b[8]), .CI(b[6]), .CO(n172), .S(n173) );
  ADDFXL U121 ( .A(b[3]), .B(b[6]), .CI(b[4]), .CO(n176), .S(n177) );
  ADDFXL U129 ( .A(n161), .B(n162), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U130 ( .A(n157), .B(n158), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U131 ( .A(n153), .B(n154), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U132 ( .A(n149), .B(n150), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U133 ( .A(n139), .B(n140), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U134 ( .A(n141), .B(n142), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U135 ( .A(n143), .B(n144), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U136 ( .A(n145), .B(n146), .CI(n43), .CO(n42), .S(product[22]) );
  ADDHXL U137 ( .A(b[3]), .B(\b[1] ), .CO(n182), .S(n183) );
  ADDFXL U138 ( .A(n165), .B(n166), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U139 ( .A(n169), .B(n170), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U140 ( .A(n173), .B(n174), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U141 ( .A(b[2]), .B(b[5]), .CI(b[3]), .CO(n178), .S(n179) );
  ADDFXL U142 ( .A(n62), .B(\b[0] ), .CI(n183), .CO(n61), .S(product[3]) );
  ADDFXL U143 ( .A(n103), .B(n104), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U144 ( .A(n107), .B(n108), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U145 ( .A(n137), .B(n138), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U146 ( .A(n75), .B(n76), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U147 ( .A(\b[1] ), .B(b[4]), .CI(b[2]), .CO(n180), .S(n181) );
  ADDHX1 U148 ( .A(\b[0] ), .B(b[2]), .CO(n62), .S(product[2]) );
  ADDFX2 U149 ( .A(n177), .B(n178), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFX2 U150 ( .A(n181), .B(n182), .CI(n61), .CO(n60), .S(product[4]) );
  ADDFXL U151 ( .A(n135), .B(n136), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U152 ( .A(n133), .B(n134), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U153 ( .A(n131), .B(n132), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U154 ( .A(n129), .B(n130), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U155 ( .A(n127), .B(n128), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U156 ( .A(n125), .B(n126), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U157 ( .A(n123), .B(n124), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U158 ( .A(n121), .B(n122), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U159 ( .A(n119), .B(n120), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U160 ( .A(n117), .B(n118), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U161 ( .A(n115), .B(n116), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U162 ( .A(n113), .B(n114), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U163 ( .A(n111), .B(n112), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U164 ( .A(n109), .B(n110), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U165 ( .A(n101), .B(n102), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U166 ( .A(n105), .B(n106), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U167 ( .A(n85), .B(n86), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U168 ( .A(n89), .B(n90), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U169 ( .A(n93), .B(n94), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U170 ( .A(n97), .B(n98), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U171 ( .A(n77), .B(n78), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U172 ( .A(n79), .B(n80), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U173 ( .A(n81), .B(n82), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U174 ( .A(n71), .B(n72), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U175 ( .A(n73), .B(n74), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U176 ( .A(n65), .B(n66), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U177 ( .A(b[4]), .B(b[7]), .CI(b[5]), .CO(n174), .S(n175) );
  ADDFXL U178 ( .A(n167), .B(n168), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U179 ( .A(n147), .B(n148), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U180 ( .A(n87), .B(n88), .CI(n14), .CO(n13), .S(product[51]) );
  XOR2X1 U181 ( .A(n321), .B(n322), .Y(product[63]) );
  XOR2X1 U182 ( .A(n323), .B(b[63]), .Y(n321) );
  XNOR2X1 U183 ( .A(n64), .B(n2), .Y(n323) );
  XNOR2X1 U184 ( .A(b[61]), .B(b[60]), .Y(n322) );
endmodule


module GSIM_DW_mult_tc_7 ( a, b, product );
  input [4:0] a;
  input [63:0] b;
  output [68:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, \b[0] , \b[1] , n321, n322, n323;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[1] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U3 ( .A(n65), .B(n66), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U5 ( .A(n69), .B(n70), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U8 ( .A(n75), .B(n76), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U10 ( .A(n79), .B(n80), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U14 ( .A(n87), .B(n88), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U16 ( .A(n91), .B(n92), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U18 ( .A(n95), .B(n96), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U20 ( .A(n99), .B(n100), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U47 ( .A(n153), .B(n154), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U49 ( .A(n157), .B(n158), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U51 ( .A(n161), .B(n162), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U53 ( .A(n165), .B(n166), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U55 ( .A(n169), .B(n170), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U57 ( .A(n173), .B(n174), .CI(n57), .CO(n56), .S(product[8]) );
  ADDHXL U63 ( .A(\b[0] ), .B(b[2]), .CO(n62), .S(product[2]) );
  ADDFXL U65 ( .A(b[59]), .B(b[62]), .CI(b[60]), .CO(n64), .S(n65) );
  ADDFXL U66 ( .A(b[58]), .B(b[61]), .CI(b[59]), .CO(n66), .S(n67) );
  ADDFXL U67 ( .A(b[57]), .B(b[60]), .CI(b[58]), .CO(n68), .S(n69) );
  ADDFXL U68 ( .A(b[56]), .B(b[59]), .CI(b[57]), .CO(n70), .S(n71) );
  ADDFXL U69 ( .A(b[55]), .B(b[58]), .CI(b[56]), .CO(n72), .S(n73) );
  ADDFXL U70 ( .A(b[54]), .B(b[57]), .CI(b[55]), .CO(n74), .S(n75) );
  ADDFXL U71 ( .A(b[53]), .B(b[56]), .CI(b[54]), .CO(n76), .S(n77) );
  ADDFXL U72 ( .A(b[52]), .B(b[55]), .CI(b[53]), .CO(n78), .S(n79) );
  ADDFXL U73 ( .A(b[51]), .B(b[54]), .CI(b[52]), .CO(n80), .S(n81) );
  ADDFXL U74 ( .A(b[50]), .B(b[53]), .CI(b[51]), .CO(n82), .S(n83) );
  ADDFXL U75 ( .A(b[49]), .B(b[52]), .CI(b[50]), .CO(n84), .S(n85) );
  ADDFXL U76 ( .A(b[48]), .B(b[51]), .CI(b[49]), .CO(n86), .S(n87) );
  ADDFXL U77 ( .A(b[47]), .B(b[50]), .CI(b[48]), .CO(n88), .S(n89) );
  ADDFXL U78 ( .A(b[46]), .B(b[49]), .CI(b[47]), .CO(n90), .S(n91) );
  ADDFXL U79 ( .A(b[45]), .B(b[48]), .CI(b[46]), .CO(n92), .S(n93) );
  ADDFXL U80 ( .A(b[44]), .B(b[47]), .CI(b[45]), .CO(n94), .S(n95) );
  ADDFXL U81 ( .A(b[43]), .B(b[46]), .CI(b[44]), .CO(n96), .S(n97) );
  ADDFXL U82 ( .A(b[42]), .B(b[45]), .CI(b[43]), .CO(n98), .S(n99) );
  ADDFXL U83 ( .A(b[41]), .B(b[44]), .CI(b[42]), .CO(n100), .S(n101) );
  ADDFXL U84 ( .A(b[40]), .B(b[43]), .CI(b[41]), .CO(n102), .S(n103) );
  ADDFXL U85 ( .A(b[39]), .B(b[42]), .CI(b[40]), .CO(n104), .S(n105) );
  ADDFXL U86 ( .A(b[38]), .B(b[41]), .CI(b[39]), .CO(n106), .S(n107) );
  ADDFXL U87 ( .A(b[37]), .B(b[40]), .CI(b[38]), .CO(n108), .S(n109) );
  ADDFXL U88 ( .A(b[36]), .B(b[39]), .CI(b[37]), .CO(n110), .S(n111) );
  ADDFXL U89 ( .A(b[35]), .B(b[38]), .CI(b[36]), .CO(n112), .S(n113) );
  ADDFXL U90 ( .A(b[34]), .B(b[37]), .CI(b[35]), .CO(n114), .S(n115) );
  ADDFXL U91 ( .A(b[33]), .B(b[36]), .CI(b[34]), .CO(n116), .S(n117) );
  ADDFXL U92 ( .A(b[32]), .B(b[35]), .CI(b[33]), .CO(n118), .S(n119) );
  ADDFXL U93 ( .A(b[31]), .B(b[34]), .CI(b[32]), .CO(n120), .S(n121) );
  ADDFXL U94 ( .A(b[30]), .B(b[33]), .CI(b[31]), .CO(n122), .S(n123) );
  ADDFXL U95 ( .A(b[29]), .B(b[32]), .CI(b[30]), .CO(n124), .S(n125) );
  ADDFXL U96 ( .A(b[28]), .B(b[31]), .CI(b[29]), .CO(n126), .S(n127) );
  ADDFXL U97 ( .A(b[27]), .B(b[30]), .CI(b[28]), .CO(n128), .S(n129) );
  ADDFXL U98 ( .A(b[26]), .B(b[29]), .CI(b[27]), .CO(n130), .S(n131) );
  ADDFXL U99 ( .A(b[25]), .B(b[28]), .CI(b[26]), .CO(n132), .S(n133) );
  ADDFXL U100 ( .A(b[24]), .B(b[27]), .CI(b[25]), .CO(n134), .S(n135) );
  ADDFXL U101 ( .A(b[23]), .B(b[26]), .CI(b[24]), .CO(n136), .S(n137) );
  ADDFXL U102 ( .A(b[22]), .B(b[25]), .CI(b[23]), .CO(n138), .S(n139) );
  ADDFXL U103 ( .A(b[21]), .B(b[24]), .CI(b[22]), .CO(n140), .S(n141) );
  ADDFXL U104 ( .A(b[20]), .B(b[23]), .CI(b[21]), .CO(n142), .S(n143) );
  ADDFXL U105 ( .A(b[19]), .B(b[22]), .CI(b[20]), .CO(n144), .S(n145) );
  ADDFXL U106 ( .A(b[18]), .B(b[21]), .CI(b[19]), .CO(n146), .S(n147) );
  ADDFXL U107 ( .A(b[17]), .B(b[20]), .CI(b[18]), .CO(n148), .S(n149) );
  ADDFXL U108 ( .A(b[16]), .B(b[19]), .CI(b[17]), .CO(n150), .S(n151) );
  ADDFXL U109 ( .A(b[15]), .B(b[18]), .CI(b[16]), .CO(n152), .S(n153) );
  ADDFXL U110 ( .A(b[14]), .B(b[17]), .CI(b[15]), .CO(n154), .S(n155) );
  ADDFXL U111 ( .A(b[13]), .B(b[16]), .CI(b[14]), .CO(n156), .S(n157) );
  ADDFXL U112 ( .A(b[12]), .B(b[15]), .CI(b[13]), .CO(n158), .S(n159) );
  ADDFXL U113 ( .A(b[11]), .B(b[14]), .CI(b[12]), .CO(n160), .S(n161) );
  ADDFXL U114 ( .A(b[10]), .B(b[13]), .CI(b[11]), .CO(n162), .S(n163) );
  ADDFXL U115 ( .A(b[9]), .B(b[12]), .CI(b[10]), .CO(n164), .S(n165) );
  ADDFXL U116 ( .A(b[8]), .B(b[11]), .CI(b[9]), .CO(n166), .S(n167) );
  ADDFXL U117 ( .A(b[7]), .B(b[10]), .CI(b[8]), .CO(n168), .S(n169) );
  ADDFXL U118 ( .A(b[6]), .B(b[9]), .CI(b[7]), .CO(n170), .S(n171) );
  ADDFXL U119 ( .A(b[5]), .B(b[8]), .CI(b[6]), .CO(n172), .S(n173) );
  ADDFXL U120 ( .A(b[4]), .B(b[7]), .CI(b[5]), .CO(n174), .S(n175) );
  ADDFXL U121 ( .A(b[3]), .B(b[6]), .CI(b[4]), .CO(n176), .S(n177) );
  ADDFXL U123 ( .A(\b[1] ), .B(b[4]), .CI(b[2]), .CO(n180), .S(n181) );
  ADDHXL U124 ( .A(b[3]), .B(\b[1] ), .CO(n182), .S(n183) );
  ADDFXL U129 ( .A(b[2]), .B(b[5]), .CI(b[3]), .CO(n178), .S(n179) );
  ADDFXL U130 ( .A(n159), .B(n160), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U131 ( .A(n155), .B(n156), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U132 ( .A(n151), .B(n152), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U133 ( .A(n181), .B(n182), .CI(n61), .CO(n60), .S(product[4]) );
  ADDFXL U134 ( .A(n163), .B(n164), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U135 ( .A(n171), .B(n172), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U136 ( .A(n167), .B(n168), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U137 ( .A(n175), .B(n176), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U138 ( .A(n62), .B(\b[0] ), .CI(n183), .CO(n61), .S(product[3]) );
  ADDFXL U139 ( .A(n149), .B(n150), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U140 ( .A(n145), .B(n146), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U141 ( .A(n141), .B(n142), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U142 ( .A(n137), .B(n138), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U143 ( .A(n133), .B(n134), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U144 ( .A(n129), .B(n130), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U145 ( .A(n125), .B(n126), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U146 ( .A(n121), .B(n122), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U147 ( .A(n117), .B(n118), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U148 ( .A(n113), .B(n114), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U149 ( .A(n109), .B(n110), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U150 ( .A(n105), .B(n106), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U151 ( .A(n101), .B(n102), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U152 ( .A(n97), .B(n98), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U153 ( .A(n93), .B(n94), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U154 ( .A(n89), .B(n90), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U155 ( .A(n85), .B(n86), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U156 ( .A(n81), .B(n82), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U157 ( .A(n73), .B(n74), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U158 ( .A(n67), .B(n68), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U159 ( .A(n77), .B(n78), .CI(n9), .CO(n8), .S(product[56]) );
  XNOR2XL U160 ( .A(b[61]), .B(b[60]), .Y(n322) );
  ADDFXL U161 ( .A(n147), .B(n148), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U162 ( .A(n143), .B(n144), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U163 ( .A(n139), .B(n140), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U164 ( .A(n135), .B(n136), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U165 ( .A(n131), .B(n132), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U166 ( .A(n127), .B(n128), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U167 ( .A(n123), .B(n124), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U168 ( .A(n119), .B(n120), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U169 ( .A(n115), .B(n116), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U170 ( .A(n111), .B(n112), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U171 ( .A(n107), .B(n108), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U172 ( .A(n71), .B(n72), .CI(n6), .CO(n5), .S(product[59]) );
  XOR2X1 U173 ( .A(n323), .B(b[63]), .Y(n321) );
  XNOR2X1 U174 ( .A(n64), .B(n2), .Y(n323) );
  ADDFXL U175 ( .A(n103), .B(n104), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U176 ( .A(n83), .B(n84), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U177 ( .A(n179), .B(n180), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U178 ( .A(n177), .B(n178), .CI(n59), .CO(n58), .S(product[6]) );
  XOR2X1 U179 ( .A(n321), .B(n322), .Y(product[63]) );
endmodule


module GSIM_DW_mult_tc_6 ( a, b, product );
  input [3:0] a;
  input [63:0] b;
  output [67:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, \b[0] , \b[1] , n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318;
  assign product[1] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[2] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U4 ( .A(b[60]), .B(n316), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U5 ( .A(b[59]), .B(n315), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U6 ( .A(b[58]), .B(n314), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U7 ( .A(b[57]), .B(n313), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U8 ( .A(b[56]), .B(n312), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U9 ( .A(b[55]), .B(n311), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U10 ( .A(b[54]), .B(n310), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U11 ( .A(b[53]), .B(n309), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U12 ( .A(b[52]), .B(n308), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U17 ( .A(b[47]), .B(n303), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U18 ( .A(b[46]), .B(n302), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U19 ( .A(b[45]), .B(n301), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U20 ( .A(b[44]), .B(n300), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U21 ( .A(b[43]), .B(n299), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U22 ( .A(b[42]), .B(n298), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U23 ( .A(b[41]), .B(n297), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U27 ( .A(b[37]), .B(n293), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U28 ( .A(b[36]), .B(n292), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U29 ( .A(b[35]), .B(n291), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U30 ( .A(b[34]), .B(n290), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U31 ( .A(b[33]), .B(n289), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U32 ( .A(b[32]), .B(n288), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U33 ( .A(b[31]), .B(n287), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U37 ( .A(b[27]), .B(n283), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U38 ( .A(b[26]), .B(n282), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U39 ( .A(b[25]), .B(n281), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U40 ( .A(b[24]), .B(n280), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U41 ( .A(b[23]), .B(n279), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U42 ( .A(b[22]), .B(n278), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U43 ( .A(b[21]), .B(n277), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U47 ( .A(b[17]), .B(n273), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U48 ( .A(b[16]), .B(n272), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U49 ( .A(b[15]), .B(n271), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U50 ( .A(b[14]), .B(n270), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U51 ( .A(b[13]), .B(n269), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U52 ( .A(b[12]), .B(n268), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U53 ( .A(b[11]), .B(n267), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U56 ( .A(b[8]), .B(n264), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U57 ( .A(b[7]), .B(n263), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U58 ( .A(b[6]), .B(n262), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U59 ( .A(b[5]), .B(n261), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U60 ( .A(b[4]), .B(n260), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFX2 U131 ( .A(b[39]), .B(n295), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U132 ( .A(b[49]), .B(n305), .CI(n15), .CO(n14), .S(product[50]) );
  CLKINVX1 U133 ( .A(b[2]), .Y(n260) );
  ADDFXL U134 ( .A(b[51]), .B(n307), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U135 ( .A(b[61]), .B(n317), .CI(n3), .CO(n2), .S(product[62]) );
  INVX1 U136 ( .A(\b[1] ), .Y(n259) );
  ADDFHX1 U137 ( .A(b[3]), .B(n259), .CI(n61), .CO(n60), .S(product[4]) );
  XOR2XL U138 ( .A(b[2]), .B(\b[0] ), .Y(product[3]) );
  ADDFXL U139 ( .A(b[10]), .B(n266), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U140 ( .A(b[20]), .B(n276), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFHX2 U141 ( .A(b[29]), .B(n285), .CI(n35), .CO(n34), .S(product[30]) );
  INVXL U142 ( .A(b[15]), .Y(n273) );
  INVXL U143 ( .A(b[24]), .Y(n282) );
  INVXL U144 ( .A(b[6]), .Y(n264) );
  INVXL U145 ( .A(b[10]), .Y(n268) );
  INVXL U146 ( .A(b[19]), .Y(n277) );
  INVXL U147 ( .A(b[20]), .Y(n278) );
  INVXL U148 ( .A(b[9]), .Y(n267) );
  INVXL U149 ( .A(b[3]), .Y(n261) );
  INVXL U150 ( .A(b[4]), .Y(n262) );
  INVXL U151 ( .A(b[5]), .Y(n263) );
  INVXL U152 ( .A(b[11]), .Y(n269) );
  INVXL U153 ( .A(b[12]), .Y(n270) );
  INVXL U154 ( .A(b[13]), .Y(n271) );
  INVXL U155 ( .A(b[14]), .Y(n272) );
  INVXL U156 ( .A(b[21]), .Y(n279) );
  INVXL U157 ( .A(b[22]), .Y(n280) );
  INVXL U158 ( .A(b[23]), .Y(n281) );
  ADDFXL U159 ( .A(b[9]), .B(n265), .CI(n55), .CO(n54), .S(product[10]) );
  INVXL U160 ( .A(b[7]), .Y(n265) );
  ADDFXL U161 ( .A(b[18]), .B(n274), .CI(n46), .CO(n45), .S(product[19]) );
  INVXL U162 ( .A(b[16]), .Y(n274) );
  ADDFXL U163 ( .A(b[19]), .B(n275), .CI(n45), .CO(n44), .S(product[20]) );
  INVXL U164 ( .A(b[17]), .Y(n275) );
  INVXL U165 ( .A(b[8]), .Y(n266) );
  INVXL U166 ( .A(b[18]), .Y(n276) );
  INVXL U167 ( .A(b[35]), .Y(n293) );
  INVXL U168 ( .A(b[44]), .Y(n302) );
  INVXL U169 ( .A(b[32]), .Y(n290) );
  INVXL U170 ( .A(b[25]), .Y(n283) );
  INVXL U171 ( .A(b[29]), .Y(n287) );
  INVXL U172 ( .A(b[30]), .Y(n288) );
  INVXL U173 ( .A(b[39]), .Y(n297) );
  INVXL U174 ( .A(b[40]), .Y(n298) );
  INVXL U175 ( .A(b[31]), .Y(n289) );
  INVXL U176 ( .A(b[33]), .Y(n291) );
  INVXL U177 ( .A(b[34]), .Y(n292) );
  INVXL U178 ( .A(b[41]), .Y(n299) );
  INVXL U179 ( .A(b[42]), .Y(n300) );
  INVXL U180 ( .A(b[43]), .Y(n301) );
  ADDFXL U181 ( .A(b[28]), .B(n284), .CI(n36), .CO(n35), .S(product[29]) );
  INVXL U182 ( .A(b[26]), .Y(n284) );
  ADDFXL U183 ( .A(b[38]), .B(n294), .CI(n26), .CO(n25), .S(product[39]) );
  INVXL U184 ( .A(b[36]), .Y(n294) );
  INVXL U185 ( .A(b[27]), .Y(n285) );
  INVXL U186 ( .A(b[37]), .Y(n295) );
  ADDFXL U187 ( .A(b[30]), .B(n286), .CI(n34), .CO(n33), .S(product[31]) );
  INVXL U188 ( .A(b[28]), .Y(n286) );
  ADDFXL U189 ( .A(b[40]), .B(n296), .CI(n24), .CO(n23), .S(product[41]) );
  INVXL U190 ( .A(b[38]), .Y(n296) );
  INVXL U191 ( .A(b[45]), .Y(n303) );
  INVXL U192 ( .A(b[58]), .Y(n316) );
  INVXL U193 ( .A(b[50]), .Y(n308) );
  INVXL U194 ( .A(b[51]), .Y(n309) );
  INVXL U195 ( .A(b[52]), .Y(n310) );
  INVXL U196 ( .A(b[53]), .Y(n311) );
  INVXL U197 ( .A(b[54]), .Y(n312) );
  INVXL U198 ( .A(b[55]), .Y(n313) );
  INVXL U199 ( .A(b[56]), .Y(n314) );
  INVXL U200 ( .A(b[57]), .Y(n315) );
  ADDFXL U201 ( .A(b[48]), .B(n304), .CI(n16), .CO(n15), .S(product[49]) );
  INVXL U202 ( .A(b[46]), .Y(n304) );
  INVXL U203 ( .A(b[59]), .Y(n317) );
  INVXL U204 ( .A(b[47]), .Y(n305) );
  ADDFXL U205 ( .A(b[50]), .B(n306), .CI(n14), .CO(n13), .S(product[51]) );
  INVXL U206 ( .A(b[48]), .Y(n306) );
  INVXL U207 ( .A(b[49]), .Y(n307) );
  XOR2XL U208 ( .A(n318), .B(b[60]), .Y(product[63]) );
  XNOR2X1 U209 ( .A(n2), .B(b[62]), .Y(n318) );
  NAND2X1 U210 ( .A(\b[0] ), .B(n260), .Y(n61) );
endmodule


module GSIM_DW01_add_483 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;
  assign SUM[15] = B[15];
  assign SUM[14] = B[14];
  assign SUM[13] = B[13];
  assign SUM[12] = B[12];
  assign SUM[11] = B[11];
  assign SUM[10] = B[10];
  assign SUM[9] = B[9];
  assign SUM[8] = B[8];
  assign SUM[7] = B[7];
  assign SUM[6] = B[6];
  assign SUM[5] = B[5];
  assign SUM[4] = B[4];
  assign SUM[3] = B[3];
  assign SUM[2] = B[2];
  assign SUM[1] = B[1];

  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(n1), .CO(carry[18]), .S(SUM[17]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  AND2X2 U1 ( .A(B[16]), .B(A[16]), .Y(n1) );
  XOR2XL U2 ( .A(B[16]), .B(A[16]), .Y(SUM[16]) );
endmodule


module GSIM_DW01_add_482 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;
  assign SUM[0] = B[0];

  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR3X2 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CMPR32X2 U1_62 ( .A(A[62]), .B(B[62]), .C(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2XL U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module GSIM_DW01_add_481 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module GSIM_DW01_add_480 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;

  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module GSIM_DW_mult_tc_12 ( a, b, product );
  input [3:0] a;
  input [63:0] b;
  output [67:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, \b[0] , \b[1] , n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318;
  assign product[1] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[2] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U4 ( .A(b[60]), .B(n316), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U5 ( .A(b[59]), .B(n315), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U6 ( .A(b[58]), .B(n314), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U7 ( .A(b[57]), .B(n313), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U8 ( .A(b[56]), .B(n312), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U9 ( .A(b[55]), .B(n311), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U11 ( .A(b[53]), .B(n309), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U12 ( .A(b[52]), .B(n308), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U13 ( .A(b[51]), .B(n307), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U14 ( .A(b[50]), .B(n306), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U15 ( .A(b[49]), .B(n305), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U16 ( .A(b[48]), .B(n304), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U17 ( .A(b[47]), .B(n303), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U18 ( .A(b[46]), .B(n302), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U19 ( .A(b[45]), .B(n301), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U21 ( .A(b[43]), .B(n299), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U22 ( .A(b[42]), .B(n298), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U23 ( .A(b[41]), .B(n297), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U24 ( .A(b[40]), .B(n296), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U25 ( .A(b[39]), .B(n295), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U26 ( .A(b[38]), .B(n294), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U27 ( .A(b[37]), .B(n293), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U28 ( .A(b[36]), .B(n292), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U29 ( .A(b[35]), .B(n291), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U31 ( .A(b[33]), .B(n289), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U32 ( .A(b[32]), .B(n288), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U33 ( .A(b[31]), .B(n287), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U34 ( .A(b[30]), .B(n286), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U35 ( .A(b[29]), .B(n285), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U36 ( .A(b[28]), .B(n284), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U37 ( .A(b[27]), .B(n283), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U38 ( .A(b[26]), .B(n282), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U39 ( .A(b[25]), .B(n281), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U41 ( .A(b[23]), .B(n279), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U42 ( .A(b[22]), .B(n278), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U43 ( .A(b[21]), .B(n277), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U44 ( .A(b[20]), .B(n276), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U45 ( .A(b[19]), .B(n275), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U46 ( .A(b[18]), .B(n274), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U47 ( .A(b[17]), .B(n273), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U48 ( .A(b[16]), .B(n272), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U49 ( .A(b[15]), .B(n271), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U51 ( .A(b[13]), .B(n269), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U52 ( .A(b[12]), .B(n268), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U53 ( .A(b[11]), .B(n267), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U54 ( .A(b[10]), .B(n266), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U55 ( .A(b[9]), .B(n265), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U56 ( .A(b[8]), .B(n264), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U57 ( .A(b[7]), .B(n263), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U58 ( .A(b[6]), .B(n262), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U59 ( .A(b[5]), .B(n261), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U131 ( .A(b[61]), .B(n317), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U132 ( .A(b[4]), .B(n260), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U133 ( .A(b[3]), .B(n259), .CI(n61), .CO(n60), .S(product[4]) );
  NAND2XL U134 ( .A(\b[0] ), .B(n260), .Y(n61) );
  ADDFXL U135 ( .A(b[14]), .B(n270), .CI(n50), .CO(n49), .S(product[15]) );
  XOR2XL U136 ( .A(b[2]), .B(\b[0] ), .Y(product[3]) );
  INVXL U137 ( .A(b[4]), .Y(n262) );
  ADDFXL U138 ( .A(b[24]), .B(n280), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFHX2 U139 ( .A(b[44]), .B(n300), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFHX2 U140 ( .A(b[54]), .B(n310), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFHX2 U141 ( .A(b[34]), .B(n290), .CI(n30), .CO(n29), .S(product[35]) );
  INVXL U142 ( .A(b[43]), .Y(n301) );
  INVXL U143 ( .A(b[44]), .Y(n302) );
  INVXL U144 ( .A(b[40]), .Y(n298) );
  INVXL U145 ( .A(b[39]), .Y(n297) );
  INVXL U146 ( .A(b[38]), .Y(n296) );
  INVXL U147 ( .A(b[37]), .Y(n295) );
  INVXL U148 ( .A(b[36]), .Y(n294) );
  INVXL U149 ( .A(b[35]), .Y(n293) );
  INVXL U150 ( .A(b[34]), .Y(n292) );
  INVXL U151 ( .A(b[33]), .Y(n291) );
  INVXL U152 ( .A(b[30]), .Y(n288) );
  INVXL U153 ( .A(b[29]), .Y(n287) );
  INVXL U154 ( .A(b[28]), .Y(n286) );
  INVXL U155 ( .A(b[13]), .Y(n271) );
  INVXL U156 ( .A(b[27]), .Y(n285) );
  INVXL U157 ( .A(b[26]), .Y(n284) );
  INVXL U158 ( .A(b[25]), .Y(n283) );
  INVXL U159 ( .A(b[24]), .Y(n282) );
  INVXL U160 ( .A(b[23]), .Y(n281) );
  INVXL U161 ( .A(b[14]), .Y(n272) );
  INVXL U162 ( .A(b[15]), .Y(n273) );
  INVXL U163 ( .A(b[16]), .Y(n274) );
  INVXL U164 ( .A(b[17]), .Y(n275) );
  INVXL U165 ( .A(b[18]), .Y(n276) );
  INVXL U166 ( .A(b[19]), .Y(n277) );
  INVXL U167 ( .A(b[20]), .Y(n278) );
  INVXL U168 ( .A(b[3]), .Y(n261) );
  INVXL U169 ( .A(b[5]), .Y(n263) );
  INVXL U170 ( .A(b[6]), .Y(n264) );
  INVXL U171 ( .A(b[7]), .Y(n265) );
  INVXL U172 ( .A(b[8]), .Y(n266) );
  INVXL U173 ( .A(b[9]), .Y(n267) );
  INVXL U174 ( .A(b[10]), .Y(n268) );
  CLKINVX1 U175 ( .A(b[58]), .Y(n316) );
  CLKINVX1 U176 ( .A(b[54]), .Y(n312) );
  CLKINVX1 U177 ( .A(b[45]), .Y(n303) );
  CLKINVX1 U178 ( .A(b[46]), .Y(n304) );
  CLKINVX1 U179 ( .A(b[47]), .Y(n305) );
  CLKINVX1 U180 ( .A(b[48]), .Y(n306) );
  CLKINVX1 U181 ( .A(b[49]), .Y(n307) );
  CLKINVX1 U182 ( .A(b[50]), .Y(n308) );
  CLKINVX1 U183 ( .A(b[53]), .Y(n311) );
  CLKINVX1 U184 ( .A(b[55]), .Y(n313) );
  CLKINVX1 U185 ( .A(b[56]), .Y(n314) );
  CLKINVX1 U186 ( .A(b[57]), .Y(n315) );
  INVXL U187 ( .A(b[11]), .Y(n269) );
  INVXL U188 ( .A(b[21]), .Y(n279) );
  INVXL U189 ( .A(b[31]), .Y(n289) );
  INVXL U190 ( .A(b[41]), .Y(n299) );
  INVXL U191 ( .A(b[51]), .Y(n309) );
  INVXL U192 ( .A(b[12]), .Y(n270) );
  INVXL U193 ( .A(b[22]), .Y(n280) );
  INVXL U194 ( .A(b[32]), .Y(n290) );
  INVXL U195 ( .A(b[42]), .Y(n300) );
  INVXL U196 ( .A(b[52]), .Y(n310) );
  INVXL U197 ( .A(b[59]), .Y(n317) );
  INVXL U198 ( .A(b[2]), .Y(n260) );
  INVX1 U199 ( .A(\b[1] ), .Y(n259) );
  XOR2X1 U200 ( .A(n318), .B(b[60]), .Y(product[63]) );
  XNOR2X1 U201 ( .A(n2), .B(b[62]), .Y(n318) );
endmodule


module GSIM_DW01_add_488 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;
  assign SUM[15] = B[15];
  assign SUM[14] = B[14];
  assign SUM[13] = B[13];
  assign SUM[12] = B[12];
  assign SUM[11] = B[11];
  assign SUM[10] = B[10];
  assign SUM[9] = B[9];
  assign SUM[8] = B[8];
  assign SUM[7] = B[7];
  assign SUM[6] = B[6];
  assign SUM[5] = B[5];
  assign SUM[4] = B[4];
  assign SUM[3] = B[3];
  assign SUM[2] = B[2];
  assign SUM[1] = B[1];

  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(n1), .CO(carry[18]), .S(SUM[17]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  AND2X2 U1 ( .A(B[16]), .B(A[16]), .Y(n1) );
  XOR2X1 U2 ( .A(B[16]), .B(A[16]), .Y(SUM[16]) );
endmodule


module GSIM_DW_mult_tc_11 ( a, b, product );
  input [3:0] a;
  input [63:0] b;
  output [67:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, \b[0] , \b[1] , n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318;
  assign product[1] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[2] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U3 ( .A(b[61]), .B(n317), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U4 ( .A(b[60]), .B(n316), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U5 ( .A(b[59]), .B(n315), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U6 ( .A(b[58]), .B(n314), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U7 ( .A(b[57]), .B(n313), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U8 ( .A(b[56]), .B(n312), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U9 ( .A(b[55]), .B(n311), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U10 ( .A(b[54]), .B(n310), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U11 ( .A(b[53]), .B(n309), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U12 ( .A(b[52]), .B(n308), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U13 ( .A(b[51]), .B(n307), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U14 ( .A(b[50]), .B(n306), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U15 ( .A(b[49]), .B(n305), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U16 ( .A(b[48]), .B(n304), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U17 ( .A(b[47]), .B(n303), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U18 ( .A(b[46]), .B(n302), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U19 ( .A(b[45]), .B(n301), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U20 ( .A(b[44]), .B(n300), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U21 ( .A(b[43]), .B(n299), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U22 ( .A(b[42]), .B(n298), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U23 ( .A(b[41]), .B(n297), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U24 ( .A(b[40]), .B(n296), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U25 ( .A(b[39]), .B(n295), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U26 ( .A(b[38]), .B(n294), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U27 ( .A(b[37]), .B(n293), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U28 ( .A(b[36]), .B(n292), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U29 ( .A(b[35]), .B(n291), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U30 ( .A(b[34]), .B(n290), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U31 ( .A(b[33]), .B(n289), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U32 ( .A(b[32]), .B(n288), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U33 ( .A(b[31]), .B(n287), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U34 ( .A(b[30]), .B(n286), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U35 ( .A(b[29]), .B(n285), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U36 ( .A(b[28]), .B(n284), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U37 ( .A(b[27]), .B(n283), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U38 ( .A(b[26]), .B(n282), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U39 ( .A(b[25]), .B(n281), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U40 ( .A(b[24]), .B(n280), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U41 ( .A(b[23]), .B(n279), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U42 ( .A(b[22]), .B(n278), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U43 ( .A(b[21]), .B(n277), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U44 ( .A(b[20]), .B(n276), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U45 ( .A(b[19]), .B(n275), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U46 ( .A(b[18]), .B(n274), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U47 ( .A(b[17]), .B(n273), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U48 ( .A(b[16]), .B(n272), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U49 ( .A(b[15]), .B(n271), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U50 ( .A(b[14]), .B(n270), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U51 ( .A(b[13]), .B(n269), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U52 ( .A(b[12]), .B(n268), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U53 ( .A(b[11]), .B(n267), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U54 ( .A(b[10]), .B(n266), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U55 ( .A(b[9]), .B(n265), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U56 ( .A(b[8]), .B(n264), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U57 ( .A(b[7]), .B(n263), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U58 ( .A(b[6]), .B(n262), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U59 ( .A(b[5]), .B(n261), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U60 ( .A(b[4]), .B(n260), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U61 ( .A(b[3]), .B(n259), .CI(n61), .CO(n60), .S(product[4]) );
  NAND2X1 U131 ( .A(\b[0] ), .B(n260), .Y(n61) );
  INVXL U132 ( .A(b[41]), .Y(n299) );
  INVXL U133 ( .A(b[42]), .Y(n300) );
  INVXL U134 ( .A(b[40]), .Y(n298) );
  INVXL U135 ( .A(b[43]), .Y(n301) );
  INVXL U136 ( .A(b[39]), .Y(n297) );
  INVXL U137 ( .A(b[38]), .Y(n296) );
  INVXL U138 ( .A(b[37]), .Y(n295) );
  INVXL U139 ( .A(b[36]), .Y(n294) );
  INVXL U140 ( .A(b[35]), .Y(n293) );
  INVXL U141 ( .A(b[34]), .Y(n292) );
  INVXL U142 ( .A(b[33]), .Y(n291) );
  INVXL U143 ( .A(b[32]), .Y(n290) );
  INVXL U144 ( .A(b[31]), .Y(n289) );
  INVXL U145 ( .A(b[30]), .Y(n288) );
  INVXL U146 ( .A(b[29]), .Y(n287) );
  INVXL U147 ( .A(b[28]), .Y(n286) );
  INVXL U148 ( .A(b[27]), .Y(n285) );
  INVXL U149 ( .A(b[26]), .Y(n284) );
  INVXL U150 ( .A(b[25]), .Y(n283) );
  INVXL U151 ( .A(b[24]), .Y(n282) );
  INVXL U152 ( .A(b[23]), .Y(n281) );
  INVXL U153 ( .A(b[22]), .Y(n280) );
  INVXL U154 ( .A(b[21]), .Y(n279) );
  INVXL U155 ( .A(b[20]), .Y(n278) );
  INVXL U156 ( .A(b[3]), .Y(n261) );
  INVXL U157 ( .A(b[4]), .Y(n262) );
  INVXL U158 ( .A(b[5]), .Y(n263) );
  INVXL U159 ( .A(b[6]), .Y(n264) );
  INVXL U160 ( .A(b[7]), .Y(n265) );
  INVXL U161 ( .A(b[8]), .Y(n266) );
  INVXL U162 ( .A(b[9]), .Y(n267) );
  INVXL U163 ( .A(b[10]), .Y(n268) );
  INVXL U164 ( .A(b[11]), .Y(n269) );
  INVXL U165 ( .A(b[12]), .Y(n270) );
  INVXL U166 ( .A(b[13]), .Y(n271) );
  INVXL U167 ( .A(b[14]), .Y(n272) );
  INVXL U168 ( .A(b[15]), .Y(n273) );
  INVXL U169 ( .A(b[16]), .Y(n274) );
  INVXL U170 ( .A(b[17]), .Y(n275) );
  INVXL U171 ( .A(b[18]), .Y(n276) );
  INVXL U172 ( .A(b[19]), .Y(n277) );
  XOR2XL U173 ( .A(b[2]), .B(\b[0] ), .Y(product[3]) );
  INVXL U174 ( .A(\b[1] ), .Y(n259) );
  CLKINVX1 U175 ( .A(b[48]), .Y(n306) );
  CLKINVX1 U176 ( .A(b[47]), .Y(n305) );
  CLKINVX1 U177 ( .A(b[49]), .Y(n307) );
  CLKINVX1 U178 ( .A(b[50]), .Y(n308) );
  CLKINVX1 U179 ( .A(b[51]), .Y(n309) );
  CLKINVX1 U180 ( .A(b[46]), .Y(n304) );
  CLKINVX1 U181 ( .A(b[44]), .Y(n302) );
  CLKINVX1 U182 ( .A(b[45]), .Y(n303) );
  CLKINVX1 U183 ( .A(b[52]), .Y(n310) );
  CLKINVX1 U184 ( .A(b[53]), .Y(n311) );
  CLKINVX1 U185 ( .A(b[54]), .Y(n312) );
  CLKINVX1 U186 ( .A(b[55]), .Y(n313) );
  CLKINVX1 U187 ( .A(b[56]), .Y(n314) );
  CLKINVX1 U188 ( .A(b[57]), .Y(n315) );
  CLKINVX1 U189 ( .A(b[58]), .Y(n316) );
  CLKINVX1 U190 ( .A(b[59]), .Y(n317) );
  INVXL U191 ( .A(b[2]), .Y(n260) );
  XOR2X1 U192 ( .A(n318), .B(b[60]), .Y(product[63]) );
  XNOR2X1 U193 ( .A(n2), .B(b[62]), .Y(n318) );
endmodule


module GSIM_DW01_add_487 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;

  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFX2 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFX2 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2XL U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module GSIM_DW_mult_tc_10 ( a, b, product );
  input [4:0] a;
  input [63:0] b;
  output [68:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, \b[0] , \b[1] , n321, n322, n323;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[1] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U3 ( .A(n65), .B(n66), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U4 ( .A(n67), .B(n68), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U6 ( .A(n71), .B(n72), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U12 ( .A(n83), .B(n84), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U14 ( .A(n87), .B(n88), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U16 ( .A(n91), .B(n92), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U18 ( .A(n95), .B(n96), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U44 ( .A(n147), .B(n148), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U46 ( .A(n151), .B(n152), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U48 ( .A(n155), .B(n156), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U52 ( .A(n163), .B(n164), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U54 ( .A(n167), .B(n168), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U56 ( .A(n171), .B(n172), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U58 ( .A(n175), .B(n176), .CI(n58), .CO(n57), .S(product[7]) );
  ADDHXL U63 ( .A(\b[0] ), .B(b[2]), .CO(n62), .S(product[2]) );
  ADDFXL U65 ( .A(b[59]), .B(b[62]), .CI(b[60]), .CO(n64), .S(n65) );
  ADDFXL U66 ( .A(b[58]), .B(b[61]), .CI(b[59]), .CO(n66), .S(n67) );
  ADDFXL U67 ( .A(b[57]), .B(b[60]), .CI(b[58]), .CO(n68), .S(n69) );
  ADDFXL U68 ( .A(b[56]), .B(b[59]), .CI(b[57]), .CO(n70), .S(n71) );
  ADDFXL U69 ( .A(b[55]), .B(b[58]), .CI(b[56]), .CO(n72), .S(n73) );
  ADDFXL U70 ( .A(b[54]), .B(b[57]), .CI(b[55]), .CO(n74), .S(n75) );
  ADDFXL U71 ( .A(b[53]), .B(b[56]), .CI(b[54]), .CO(n76), .S(n77) );
  ADDFXL U72 ( .A(b[52]), .B(b[55]), .CI(b[53]), .CO(n78), .S(n79) );
  ADDFXL U73 ( .A(b[51]), .B(b[54]), .CI(b[52]), .CO(n80), .S(n81) );
  ADDFXL U74 ( .A(b[50]), .B(b[53]), .CI(b[51]), .CO(n82), .S(n83) );
  ADDFXL U75 ( .A(b[49]), .B(b[52]), .CI(b[50]), .CO(n84), .S(n85) );
  ADDFXL U76 ( .A(b[48]), .B(b[51]), .CI(b[49]), .CO(n86), .S(n87) );
  ADDFXL U77 ( .A(b[47]), .B(b[50]), .CI(b[48]), .CO(n88), .S(n89) );
  ADDFXL U78 ( .A(b[46]), .B(b[49]), .CI(b[47]), .CO(n90), .S(n91) );
  ADDFXL U79 ( .A(b[45]), .B(b[48]), .CI(b[46]), .CO(n92), .S(n93) );
  ADDFXL U80 ( .A(b[44]), .B(b[47]), .CI(b[45]), .CO(n94), .S(n95) );
  ADDFXL U81 ( .A(b[43]), .B(b[46]), .CI(b[44]), .CO(n96), .S(n97) );
  ADDFXL U82 ( .A(b[42]), .B(b[45]), .CI(b[43]), .CO(n98), .S(n99) );
  ADDFXL U83 ( .A(b[41]), .B(b[44]), .CI(b[42]), .CO(n100), .S(n101) );
  ADDFXL U84 ( .A(b[40]), .B(b[43]), .CI(b[41]), .CO(n102), .S(n103) );
  ADDFXL U85 ( .A(b[39]), .B(b[42]), .CI(b[40]), .CO(n104), .S(n105) );
  ADDFXL U86 ( .A(b[38]), .B(b[41]), .CI(b[39]), .CO(n106), .S(n107) );
  ADDFXL U87 ( .A(b[37]), .B(b[40]), .CI(b[38]), .CO(n108), .S(n109) );
  ADDFXL U88 ( .A(b[36]), .B(b[39]), .CI(b[37]), .CO(n110), .S(n111) );
  ADDFXL U89 ( .A(b[35]), .B(b[38]), .CI(b[36]), .CO(n112), .S(n113) );
  ADDFXL U90 ( .A(b[34]), .B(b[37]), .CI(b[35]), .CO(n114), .S(n115) );
  ADDFXL U91 ( .A(b[33]), .B(b[36]), .CI(b[34]), .CO(n116), .S(n117) );
  ADDFXL U92 ( .A(b[32]), .B(b[35]), .CI(b[33]), .CO(n118), .S(n119) );
  ADDFXL U93 ( .A(b[31]), .B(b[34]), .CI(b[32]), .CO(n120), .S(n121) );
  ADDFXL U94 ( .A(b[30]), .B(b[33]), .CI(b[31]), .CO(n122), .S(n123) );
  ADDFXL U95 ( .A(b[29]), .B(b[32]), .CI(b[30]), .CO(n124), .S(n125) );
  ADDFXL U96 ( .A(b[28]), .B(b[31]), .CI(b[29]), .CO(n126), .S(n127) );
  ADDFXL U97 ( .A(b[27]), .B(b[30]), .CI(b[28]), .CO(n128), .S(n129) );
  ADDFXL U98 ( .A(b[26]), .B(b[29]), .CI(b[27]), .CO(n130), .S(n131) );
  ADDFXL U99 ( .A(b[25]), .B(b[28]), .CI(b[26]), .CO(n132), .S(n133) );
  ADDFXL U100 ( .A(b[24]), .B(b[27]), .CI(b[25]), .CO(n134), .S(n135) );
  ADDFXL U101 ( .A(b[23]), .B(b[26]), .CI(b[24]), .CO(n136), .S(n137) );
  ADDFXL U102 ( .A(b[22]), .B(b[25]), .CI(b[23]), .CO(n138), .S(n139) );
  ADDFXL U103 ( .A(b[21]), .B(b[24]), .CI(b[22]), .CO(n140), .S(n141) );
  ADDFXL U104 ( .A(b[20]), .B(b[23]), .CI(b[21]), .CO(n142), .S(n143) );
  ADDFXL U105 ( .A(b[19]), .B(b[22]), .CI(b[20]), .CO(n144), .S(n145) );
  ADDFXL U106 ( .A(b[18]), .B(b[21]), .CI(b[19]), .CO(n146), .S(n147) );
  ADDFXL U107 ( .A(b[17]), .B(b[20]), .CI(b[18]), .CO(n148), .S(n149) );
  ADDFXL U108 ( .A(b[16]), .B(b[19]), .CI(b[17]), .CO(n150), .S(n151) );
  ADDFXL U109 ( .A(b[15]), .B(b[18]), .CI(b[16]), .CO(n152), .S(n153) );
  ADDFXL U110 ( .A(b[14]), .B(b[17]), .CI(b[15]), .CO(n154), .S(n155) );
  ADDFXL U111 ( .A(b[13]), .B(b[16]), .CI(b[14]), .CO(n156), .S(n157) );
  ADDFXL U112 ( .A(b[12]), .B(b[15]), .CI(b[13]), .CO(n158), .S(n159) );
  ADDFXL U113 ( .A(b[11]), .B(b[14]), .CI(b[12]), .CO(n160), .S(n161) );
  ADDFXL U114 ( .A(b[10]), .B(b[13]), .CI(b[11]), .CO(n162), .S(n163) );
  ADDFXL U115 ( .A(b[9]), .B(b[12]), .CI(b[10]), .CO(n164), .S(n165) );
  ADDFXL U116 ( .A(b[8]), .B(b[11]), .CI(b[9]), .CO(n166), .S(n167) );
  ADDFXL U117 ( .A(b[7]), .B(b[10]), .CI(b[8]), .CO(n168), .S(n169) );
  ADDFXL U118 ( .A(b[6]), .B(b[9]), .CI(b[7]), .CO(n170), .S(n171) );
  ADDFXL U119 ( .A(b[5]), .B(b[8]), .CI(b[6]), .CO(n172), .S(n173) );
  ADDFXL U121 ( .A(b[3]), .B(b[6]), .CI(b[4]), .CO(n176), .S(n177) );
  ADDFXL U122 ( .A(b[2]), .B(b[5]), .CI(b[3]), .CO(n178), .S(n179) );
  ADDHXL U124 ( .A(b[3]), .B(\b[1] ), .CO(n182), .S(n183) );
  ADDFXL U129 ( .A(n153), .B(n154), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U130 ( .A(n149), .B(n150), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U131 ( .A(n139), .B(n140), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U132 ( .A(n141), .B(n142), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U133 ( .A(n143), .B(n144), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U134 ( .A(n145), .B(n146), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U135 ( .A(\b[1] ), .B(b[4]), .CI(b[2]), .CO(n180), .S(n181) );
  ADDFXL U136 ( .A(n165), .B(n166), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U137 ( .A(n169), .B(n170), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U138 ( .A(n177), .B(n178), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U139 ( .A(n137), .B(n138), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U140 ( .A(n181), .B(n182), .CI(n61), .CO(n60), .S(product[4]) );
  ADDFXL U141 ( .A(n173), .B(n174), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U142 ( .A(n161), .B(n162), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U143 ( .A(n157), .B(n158), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U144 ( .A(n123), .B(n124), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U145 ( .A(n127), .B(n128), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U146 ( .A(n131), .B(n132), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U147 ( .A(n135), .B(n136), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U148 ( .A(n79), .B(n80), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U149 ( .A(n119), .B(n120), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U150 ( .A(n73), .B(n74), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U151 ( .A(n69), .B(n70), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U152 ( .A(n62), .B(\b[0] ), .CI(n183), .CO(n61), .S(product[3]) );
  ADDFXL U153 ( .A(n133), .B(n134), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U154 ( .A(n129), .B(n130), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U155 ( .A(n125), .B(n126), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U156 ( .A(n121), .B(n122), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U157 ( .A(n117), .B(n118), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U158 ( .A(n115), .B(n116), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U159 ( .A(n113), .B(n114), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U160 ( .A(n111), .B(n112), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U161 ( .A(n109), .B(n110), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U162 ( .A(n107), .B(n108), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U163 ( .A(n105), .B(n106), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U164 ( .A(n97), .B(n98), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U165 ( .A(n101), .B(n102), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U166 ( .A(n103), .B(n104), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U167 ( .A(n85), .B(n86), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U168 ( .A(n89), .B(n90), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U169 ( .A(n93), .B(n94), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U170 ( .A(n81), .B(n82), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U171 ( .A(n77), .B(n78), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U172 ( .A(n75), .B(n76), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U173 ( .A(b[4]), .B(b[7]), .CI(b[5]), .CO(n174), .S(n175) );
  ADDFXL U174 ( .A(n179), .B(n180), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U175 ( .A(n159), .B(n160), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U176 ( .A(n99), .B(n100), .CI(n20), .CO(n19), .S(product[45]) );
  XOR2X1 U177 ( .A(n321), .B(n322), .Y(product[63]) );
  XOR2X1 U178 ( .A(n323), .B(b[63]), .Y(n321) );
  XNOR2X1 U179 ( .A(n64), .B(n2), .Y(n323) );
  XNOR2X1 U180 ( .A(b[61]), .B(b[60]), .Y(n322) );
endmodule


module GSIM_DW_mult_tc_9 ( a, b, product );
  input [4:0] a;
  input [63:0] b;
  output [68:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, \b[0] , \b[1] , n321, n322, n323;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[1] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U3 ( .A(n65), .B(n66), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U15 ( .A(n89), .B(n90), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U17 ( .A(n93), .B(n94), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U19 ( .A(n97), .B(n98), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U21 ( .A(n101), .B(n102), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U47 ( .A(n153), .B(n154), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U49 ( .A(n157), .B(n158), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U51 ( .A(n161), .B(n162), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U53 ( .A(n165), .B(n166), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U55 ( .A(n169), .B(n170), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U57 ( .A(n173), .B(n174), .CI(n57), .CO(n56), .S(product[8]) );
  ADDHXL U63 ( .A(\b[0] ), .B(b[2]), .CO(n62), .S(product[2]) );
  ADDFXL U65 ( .A(b[59]), .B(b[62]), .CI(b[60]), .CO(n64), .S(n65) );
  ADDFXL U66 ( .A(b[58]), .B(b[61]), .CI(b[59]), .CO(n66), .S(n67) );
  ADDFXL U67 ( .A(b[57]), .B(b[60]), .CI(b[58]), .CO(n68), .S(n69) );
  ADDFXL U68 ( .A(b[56]), .B(b[59]), .CI(b[57]), .CO(n70), .S(n71) );
  ADDFXL U69 ( .A(b[55]), .B(b[58]), .CI(b[56]), .CO(n72), .S(n73) );
  ADDFXL U70 ( .A(b[54]), .B(b[57]), .CI(b[55]), .CO(n74), .S(n75) );
  ADDFXL U71 ( .A(b[53]), .B(b[56]), .CI(b[54]), .CO(n76), .S(n77) );
  ADDFXL U72 ( .A(b[52]), .B(b[55]), .CI(b[53]), .CO(n78), .S(n79) );
  ADDFXL U73 ( .A(b[51]), .B(b[54]), .CI(b[52]), .CO(n80), .S(n81) );
  ADDFXL U74 ( .A(b[50]), .B(b[53]), .CI(b[51]), .CO(n82), .S(n83) );
  ADDFXL U75 ( .A(b[49]), .B(b[52]), .CI(b[50]), .CO(n84), .S(n85) );
  ADDFXL U76 ( .A(b[48]), .B(b[51]), .CI(b[49]), .CO(n86), .S(n87) );
  ADDFXL U77 ( .A(b[47]), .B(b[50]), .CI(b[48]), .CO(n88), .S(n89) );
  ADDFXL U78 ( .A(b[46]), .B(b[49]), .CI(b[47]), .CO(n90), .S(n91) );
  ADDFXL U79 ( .A(b[45]), .B(b[48]), .CI(b[46]), .CO(n92), .S(n93) );
  ADDFXL U80 ( .A(b[44]), .B(b[47]), .CI(b[45]), .CO(n94), .S(n95) );
  ADDFXL U81 ( .A(b[43]), .B(b[46]), .CI(b[44]), .CO(n96), .S(n97) );
  ADDFXL U82 ( .A(b[42]), .B(b[45]), .CI(b[43]), .CO(n98), .S(n99) );
  ADDFXL U83 ( .A(b[41]), .B(b[44]), .CI(b[42]), .CO(n100), .S(n101) );
  ADDFXL U84 ( .A(b[40]), .B(b[43]), .CI(b[41]), .CO(n102), .S(n103) );
  ADDFXL U85 ( .A(b[39]), .B(b[42]), .CI(b[40]), .CO(n104), .S(n105) );
  ADDFXL U86 ( .A(b[38]), .B(b[41]), .CI(b[39]), .CO(n106), .S(n107) );
  ADDFXL U87 ( .A(b[37]), .B(b[40]), .CI(b[38]), .CO(n108), .S(n109) );
  ADDFXL U88 ( .A(b[36]), .B(b[39]), .CI(b[37]), .CO(n110), .S(n111) );
  ADDFXL U89 ( .A(b[35]), .B(b[38]), .CI(b[36]), .CO(n112), .S(n113) );
  ADDFXL U90 ( .A(b[34]), .B(b[37]), .CI(b[35]), .CO(n114), .S(n115) );
  ADDFXL U91 ( .A(b[33]), .B(b[36]), .CI(b[34]), .CO(n116), .S(n117) );
  ADDFXL U92 ( .A(b[32]), .B(b[35]), .CI(b[33]), .CO(n118), .S(n119) );
  ADDFXL U93 ( .A(b[31]), .B(b[34]), .CI(b[32]), .CO(n120), .S(n121) );
  ADDFXL U94 ( .A(b[30]), .B(b[33]), .CI(b[31]), .CO(n122), .S(n123) );
  ADDFXL U95 ( .A(b[29]), .B(b[32]), .CI(b[30]), .CO(n124), .S(n125) );
  ADDFXL U96 ( .A(b[28]), .B(b[31]), .CI(b[29]), .CO(n126), .S(n127) );
  ADDFXL U97 ( .A(b[27]), .B(b[30]), .CI(b[28]), .CO(n128), .S(n129) );
  ADDFXL U98 ( .A(b[26]), .B(b[29]), .CI(b[27]), .CO(n130), .S(n131) );
  ADDFXL U99 ( .A(b[25]), .B(b[28]), .CI(b[26]), .CO(n132), .S(n133) );
  ADDFXL U100 ( .A(b[24]), .B(b[27]), .CI(b[25]), .CO(n134), .S(n135) );
  ADDFXL U101 ( .A(b[23]), .B(b[26]), .CI(b[24]), .CO(n136), .S(n137) );
  ADDFXL U102 ( .A(b[22]), .B(b[25]), .CI(b[23]), .CO(n138), .S(n139) );
  ADDFXL U103 ( .A(b[21]), .B(b[24]), .CI(b[22]), .CO(n140), .S(n141) );
  ADDFXL U104 ( .A(b[20]), .B(b[23]), .CI(b[21]), .CO(n142), .S(n143) );
  ADDFXL U105 ( .A(b[19]), .B(b[22]), .CI(b[20]), .CO(n144), .S(n145) );
  ADDFXL U106 ( .A(b[18]), .B(b[21]), .CI(b[19]), .CO(n146), .S(n147) );
  ADDFXL U107 ( .A(b[17]), .B(b[20]), .CI(b[18]), .CO(n148), .S(n149) );
  ADDFXL U108 ( .A(b[16]), .B(b[19]), .CI(b[17]), .CO(n150), .S(n151) );
  ADDFXL U109 ( .A(b[15]), .B(b[18]), .CI(b[16]), .CO(n152), .S(n153) );
  ADDFXL U110 ( .A(b[14]), .B(b[17]), .CI(b[15]), .CO(n154), .S(n155) );
  ADDFXL U111 ( .A(b[13]), .B(b[16]), .CI(b[14]), .CO(n156), .S(n157) );
  ADDFXL U112 ( .A(b[12]), .B(b[15]), .CI(b[13]), .CO(n158), .S(n159) );
  ADDFXL U113 ( .A(b[11]), .B(b[14]), .CI(b[12]), .CO(n160), .S(n161) );
  ADDFXL U114 ( .A(b[10]), .B(b[13]), .CI(b[11]), .CO(n162), .S(n163) );
  ADDFXL U115 ( .A(b[9]), .B(b[12]), .CI(b[10]), .CO(n164), .S(n165) );
  ADDFXL U116 ( .A(b[8]), .B(b[11]), .CI(b[9]), .CO(n166), .S(n167) );
  ADDFXL U117 ( .A(b[7]), .B(b[10]), .CI(b[8]), .CO(n168), .S(n169) );
  ADDFXL U118 ( .A(b[6]), .B(b[9]), .CI(b[7]), .CO(n170), .S(n171) );
  ADDFXL U119 ( .A(b[5]), .B(b[8]), .CI(b[6]), .CO(n172), .S(n173) );
  ADDFXL U120 ( .A(b[4]), .B(b[7]), .CI(b[5]), .CO(n174), .S(n175) );
  ADDFXL U121 ( .A(b[3]), .B(b[6]), .CI(b[4]), .CO(n176), .S(n177) );
  ADDFXL U123 ( .A(\b[1] ), .B(b[4]), .CI(b[2]), .CO(n180), .S(n181) );
  ADDHXL U124 ( .A(b[3]), .B(\b[1] ), .CO(n182), .S(n183) );
  ADDFXL U129 ( .A(b[2]), .B(b[5]), .CI(b[3]), .CO(n178), .S(n179) );
  ADDFXL U130 ( .A(n159), .B(n160), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U131 ( .A(n155), .B(n156), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U132 ( .A(n151), .B(n152), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U133 ( .A(n149), .B(n150), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U134 ( .A(n147), .B(n148), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U135 ( .A(n163), .B(n164), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U136 ( .A(n171), .B(n172), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U137 ( .A(n167), .B(n168), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U138 ( .A(n175), .B(n176), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U139 ( .A(n62), .B(\b[0] ), .CI(n183), .CO(n61), .S(product[3]) );
  ADDFXL U140 ( .A(n181), .B(n182), .CI(n61), .CO(n60), .S(product[4]) );
  ADDFXL U141 ( .A(n145), .B(n146), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U142 ( .A(n141), .B(n142), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U143 ( .A(n137), .B(n138), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U144 ( .A(n133), .B(n134), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U145 ( .A(n129), .B(n130), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U146 ( .A(n125), .B(n126), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U147 ( .A(n121), .B(n122), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U148 ( .A(n117), .B(n118), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U149 ( .A(n113), .B(n114), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U150 ( .A(n109), .B(n110), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U151 ( .A(n105), .B(n106), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U152 ( .A(n99), .B(n100), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U153 ( .A(n95), .B(n96), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U154 ( .A(n91), .B(n92), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U155 ( .A(n77), .B(n78), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U156 ( .A(n73), .B(n74), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U157 ( .A(n75), .B(n76), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U158 ( .A(n87), .B(n88), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U159 ( .A(n81), .B(n82), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U160 ( .A(n69), .B(n70), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U161 ( .A(n67), .B(n68), .CI(n4), .CO(n3), .S(product[61]) );
  XOR2X1 U162 ( .A(n323), .B(b[63]), .Y(n321) );
  XNOR2XL U163 ( .A(b[61]), .B(b[60]), .Y(n322) );
  ADDFXL U164 ( .A(n143), .B(n144), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U165 ( .A(n135), .B(n136), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U166 ( .A(n139), .B(n140), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U167 ( .A(n127), .B(n128), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U168 ( .A(n131), .B(n132), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U169 ( .A(n123), .B(n124), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U170 ( .A(n115), .B(n116), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U171 ( .A(n119), .B(n120), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U172 ( .A(n107), .B(n108), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U173 ( .A(n111), .B(n112), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U174 ( .A(n103), .B(n104), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U175 ( .A(n79), .B(n80), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U176 ( .A(n83), .B(n84), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U177 ( .A(n71), .B(n72), .CI(n6), .CO(n5), .S(product[59]) );
  XNOR2X1 U178 ( .A(n64), .B(n2), .Y(n323) );
  ADDFXL U179 ( .A(n179), .B(n180), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U180 ( .A(n177), .B(n178), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U181 ( .A(n85), .B(n86), .CI(n13), .CO(n12), .S(product[52]) );
  XOR2X1 U182 ( .A(n321), .B(n322), .Y(product[63]) );
endmodule


module GSIM_DW01_add_486 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;
  assign SUM[0] = B[0];

  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  CMPR32X2 U1_62 ( .A(A[62]), .B(B[62]), .C(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2XL U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module GSIM_DW01_add_485 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  XOR3X2 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module GSIM_DW01_add_484 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;

  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFHX2 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module GSIM_DW_mult_tc_17 ( a, b, product );
  input [3:0] a;
  input [63:0] b;
  output [67:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, \b[0] , \b[1] , n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318;
  assign product[1] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[2] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U3 ( .A(b[61]), .B(n317), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U4 ( .A(b[60]), .B(n316), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U5 ( .A(b[59]), .B(n315), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U6 ( .A(b[58]), .B(n314), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U7 ( .A(b[57]), .B(n313), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U8 ( .A(b[56]), .B(n312), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U9 ( .A(b[55]), .B(n311), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U10 ( .A(b[54]), .B(n310), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U11 ( .A(b[53]), .B(n309), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U12 ( .A(b[52]), .B(n308), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U13 ( .A(b[51]), .B(n307), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U14 ( .A(b[50]), .B(n306), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U15 ( .A(b[49]), .B(n305), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U16 ( .A(b[48]), .B(n304), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U17 ( .A(b[47]), .B(n303), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U18 ( .A(b[46]), .B(n302), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U19 ( .A(b[45]), .B(n301), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U20 ( .A(b[44]), .B(n300), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U21 ( .A(b[43]), .B(n299), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U22 ( .A(b[42]), .B(n298), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U23 ( .A(b[41]), .B(n297), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U24 ( .A(b[40]), .B(n296), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U25 ( .A(b[39]), .B(n295), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U26 ( .A(b[38]), .B(n294), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U27 ( .A(b[37]), .B(n293), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U28 ( .A(b[36]), .B(n292), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U29 ( .A(b[35]), .B(n291), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U30 ( .A(b[34]), .B(n290), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U31 ( .A(b[33]), .B(n289), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U32 ( .A(b[32]), .B(n288), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U33 ( .A(b[31]), .B(n287), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U34 ( .A(b[30]), .B(n286), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U35 ( .A(b[29]), .B(n285), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U36 ( .A(b[28]), .B(n284), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U37 ( .A(b[27]), .B(n283), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U38 ( .A(b[26]), .B(n282), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U39 ( .A(b[25]), .B(n281), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U40 ( .A(b[24]), .B(n280), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U41 ( .A(b[23]), .B(n279), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U42 ( .A(b[22]), .B(n278), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U43 ( .A(b[21]), .B(n277), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U44 ( .A(b[20]), .B(n276), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U45 ( .A(b[19]), .B(n275), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U46 ( .A(b[18]), .B(n274), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U47 ( .A(b[17]), .B(n273), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U48 ( .A(b[16]), .B(n272), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U49 ( .A(b[15]), .B(n271), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U50 ( .A(b[14]), .B(n270), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U51 ( .A(b[13]), .B(n269), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U52 ( .A(b[12]), .B(n268), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U53 ( .A(b[11]), .B(n267), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U54 ( .A(b[10]), .B(n266), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U55 ( .A(b[9]), .B(n265), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U56 ( .A(b[8]), .B(n264), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U57 ( .A(b[7]), .B(n263), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U58 ( .A(b[6]), .B(n262), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U59 ( .A(b[5]), .B(n261), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U60 ( .A(b[4]), .B(n260), .CI(n60), .CO(n59), .S(product[5]) );
  CLKINVX1 U131 ( .A(b[3]), .Y(n261) );
  ADDFXL U132 ( .A(b[3]), .B(n259), .CI(n61), .CO(n60), .S(product[4]) );
  XOR2XL U133 ( .A(b[2]), .B(\b[0] ), .Y(product[3]) );
  INVXL U134 ( .A(\b[1] ), .Y(n259) );
  NAND2XL U135 ( .A(\b[0] ), .B(n260), .Y(n61) );
  INVXL U136 ( .A(b[12]), .Y(n270) );
  INVXL U137 ( .A(b[22]), .Y(n280) );
  INVXL U138 ( .A(b[32]), .Y(n290) );
  INVXL U139 ( .A(b[42]), .Y(n300) );
  INVXL U140 ( .A(b[52]), .Y(n310) );
  INVXL U141 ( .A(b[4]), .Y(n262) );
  INVXL U142 ( .A(b[11]), .Y(n269) );
  INVXL U143 ( .A(b[21]), .Y(n279) );
  INVXL U144 ( .A(b[31]), .Y(n289) );
  INVXL U145 ( .A(b[41]), .Y(n299) );
  INVXL U146 ( .A(b[51]), .Y(n309) );
  INVXL U147 ( .A(b[14]), .Y(n272) );
  INVXL U148 ( .A(b[24]), .Y(n282) );
  INVXL U149 ( .A(b[34]), .Y(n292) );
  INVXL U150 ( .A(b[44]), .Y(n302) );
  INVXL U151 ( .A(b[54]), .Y(n312) );
  INVXL U152 ( .A(b[5]), .Y(n263) );
  INVXL U153 ( .A(b[6]), .Y(n264) );
  INVXL U154 ( .A(b[7]), .Y(n265) );
  INVXL U155 ( .A(b[8]), .Y(n266) );
  INVXL U156 ( .A(b[9]), .Y(n267) );
  INVXL U157 ( .A(b[10]), .Y(n268) );
  INVXL U158 ( .A(b[13]), .Y(n271) );
  INVXL U159 ( .A(b[15]), .Y(n273) );
  INVXL U160 ( .A(b[16]), .Y(n274) );
  INVXL U161 ( .A(b[17]), .Y(n275) );
  INVXL U162 ( .A(b[18]), .Y(n276) );
  INVXL U163 ( .A(b[19]), .Y(n277) );
  INVXL U164 ( .A(b[20]), .Y(n278) );
  INVXL U165 ( .A(b[23]), .Y(n281) );
  INVXL U166 ( .A(b[25]), .Y(n283) );
  INVXL U167 ( .A(b[26]), .Y(n284) );
  INVXL U168 ( .A(b[27]), .Y(n285) );
  INVXL U169 ( .A(b[28]), .Y(n286) );
  INVXL U170 ( .A(b[29]), .Y(n287) );
  INVXL U171 ( .A(b[30]), .Y(n288) );
  INVXL U172 ( .A(b[33]), .Y(n291) );
  INVXL U173 ( .A(b[35]), .Y(n293) );
  INVXL U174 ( .A(b[36]), .Y(n294) );
  INVXL U175 ( .A(b[37]), .Y(n295) );
  INVXL U176 ( .A(b[38]), .Y(n296) );
  INVXL U177 ( .A(b[39]), .Y(n297) );
  INVXL U178 ( .A(b[40]), .Y(n298) );
  INVXL U179 ( .A(b[43]), .Y(n301) );
  INVXL U180 ( .A(b[45]), .Y(n303) );
  INVXL U181 ( .A(b[46]), .Y(n304) );
  INVXL U182 ( .A(b[47]), .Y(n305) );
  INVXL U183 ( .A(b[48]), .Y(n306) );
  INVXL U184 ( .A(b[49]), .Y(n307) );
  INVXL U185 ( .A(b[50]), .Y(n308) );
  INVXL U186 ( .A(b[53]), .Y(n311) );
  INVXL U187 ( .A(b[55]), .Y(n313) );
  INVXL U188 ( .A(b[56]), .Y(n314) );
  INVXL U189 ( .A(b[57]), .Y(n315) );
  INVXL U190 ( .A(b[58]), .Y(n316) );
  INVXL U191 ( .A(b[59]), .Y(n317) );
  INVXL U192 ( .A(b[2]), .Y(n260) );
  XOR2X1 U193 ( .A(n318), .B(b[60]), .Y(product[63]) );
  XNOR2X1 U194 ( .A(n2), .B(b[62]), .Y(n318) );
endmodule


module GSIM_DW01_add_495 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;
  assign SUM[15] = B[15];
  assign SUM[14] = B[14];
  assign SUM[13] = B[13];
  assign SUM[12] = B[12];
  assign SUM[11] = B[11];
  assign SUM[10] = B[10];
  assign SUM[9] = B[9];
  assign SUM[8] = B[8];
  assign SUM[7] = B[7];
  assign SUM[6] = B[6];
  assign SUM[5] = B[5];
  assign SUM[4] = B[4];
  assign SUM[3] = B[3];
  assign SUM[2] = B[2];
  assign SUM[1] = B[1];

  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(n1), .CO(carry[18]), .S(SUM[17]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  AND2X2 U1 ( .A(B[16]), .B(A[16]), .Y(n1) );
  XOR2XL U2 ( .A(B[16]), .B(A[16]), .Y(SUM[16]) );
endmodule


module GSIM_DW_mult_tc_16 ( a, b, product );
  input [4:0] a;
  input [63:0] b;
  output [68:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, \b[0] , \b[1] , n321, n322, n323;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[1] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U3 ( .A(n65), .B(n66), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U13 ( .A(n85), .B(n86), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U15 ( .A(n89), .B(n90), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U17 ( .A(n93), .B(n94), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U19 ( .A(n97), .B(n98), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U21 ( .A(n101), .B(n102), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U23 ( .A(n105), .B(n106), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U25 ( .A(n109), .B(n110), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U27 ( .A(n113), .B(n114), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U29 ( .A(n117), .B(n118), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U31 ( .A(n121), .B(n122), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U50 ( .A(n159), .B(n160), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U52 ( .A(n163), .B(n164), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U54 ( .A(n167), .B(n168), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U56 ( .A(n171), .B(n172), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U58 ( .A(n175), .B(n176), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U60 ( .A(n179), .B(n180), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U62 ( .A(n62), .B(\b[0] ), .CI(n183), .CO(n61), .S(product[3]) );
  ADDHXL U63 ( .A(\b[0] ), .B(b[2]), .CO(n62), .S(product[2]) );
  ADDFXL U65 ( .A(b[59]), .B(b[62]), .CI(b[60]), .CO(n64), .S(n65) );
  ADDFXL U66 ( .A(b[58]), .B(b[61]), .CI(b[59]), .CO(n66), .S(n67) );
  ADDFXL U68 ( .A(b[56]), .B(b[59]), .CI(b[57]), .CO(n70), .S(n71) );
  ADDFXL U69 ( .A(b[55]), .B(b[58]), .CI(b[56]), .CO(n72), .S(n73) );
  ADDFXL U71 ( .A(b[53]), .B(b[56]), .CI(b[54]), .CO(n76), .S(n77) );
  ADDFXL U72 ( .A(b[52]), .B(b[55]), .CI(b[53]), .CO(n78), .S(n79) );
  ADDFXL U74 ( .A(b[50]), .B(b[53]), .CI(b[51]), .CO(n82), .S(n83) );
  ADDFXL U75 ( .A(b[49]), .B(b[52]), .CI(b[50]), .CO(n84), .S(n85) );
  ADDFXL U78 ( .A(b[46]), .B(b[49]), .CI(b[47]), .CO(n90), .S(n91) );
  ADDFXL U79 ( .A(b[45]), .B(b[48]), .CI(b[46]), .CO(n92), .S(n93) );
  ADDFXL U80 ( .A(b[44]), .B(b[47]), .CI(b[45]), .CO(n94), .S(n95) );
  ADDFXL U81 ( .A(b[43]), .B(b[46]), .CI(b[44]), .CO(n96), .S(n97) );
  ADDFXL U83 ( .A(b[41]), .B(b[44]), .CI(b[42]), .CO(n100), .S(n101) );
  ADDFXL U84 ( .A(b[40]), .B(b[43]), .CI(b[41]), .CO(n102), .S(n103) );
  ADDFXL U86 ( .A(b[38]), .B(b[41]), .CI(b[39]), .CO(n106), .S(n107) );
  ADDFXL U87 ( .A(b[37]), .B(b[40]), .CI(b[38]), .CO(n108), .S(n109) );
  ADDFXL U89 ( .A(b[35]), .B(b[38]), .CI(b[36]), .CO(n112), .S(n113) );
  ADDFXL U90 ( .A(b[34]), .B(b[37]), .CI(b[35]), .CO(n114), .S(n115) );
  ADDFXL U92 ( .A(b[32]), .B(b[35]), .CI(b[33]), .CO(n118), .S(n119) );
  ADDFXL U93 ( .A(b[31]), .B(b[34]), .CI(b[32]), .CO(n120), .S(n121) );
  ADDFXL U95 ( .A(b[29]), .B(b[32]), .CI(b[30]), .CO(n124), .S(n125) );
  ADDFXL U96 ( .A(b[28]), .B(b[31]), .CI(b[29]), .CO(n126), .S(n127) );
  ADDFXL U97 ( .A(b[27]), .B(b[30]), .CI(b[28]), .CO(n128), .S(n129) );
  ADDFXL U100 ( .A(b[24]), .B(b[27]), .CI(b[25]), .CO(n134), .S(n135) );
  ADDFXL U101 ( .A(b[23]), .B(b[26]), .CI(b[24]), .CO(n136), .S(n137) );
  ADDFXL U103 ( .A(b[21]), .B(b[24]), .CI(b[22]), .CO(n140), .S(n141) );
  ADDFXL U104 ( .A(b[20]), .B(b[23]), .CI(b[21]), .CO(n142), .S(n143) );
  ADDFXL U105 ( .A(b[19]), .B(b[22]), .CI(b[20]), .CO(n144), .S(n145) );
  ADDFXL U108 ( .A(b[16]), .B(b[19]), .CI(b[17]), .CO(n150), .S(n151) );
  ADDFXL U109 ( .A(b[15]), .B(b[18]), .CI(b[16]), .CO(n152), .S(n153) );
  ADDFXL U111 ( .A(b[13]), .B(b[16]), .CI(b[14]), .CO(n156), .S(n157) );
  ADDFXL U112 ( .A(b[12]), .B(b[15]), .CI(b[13]), .CO(n158), .S(n159) );
  ADDFXL U119 ( .A(b[5]), .B(b[8]), .CI(b[6]), .CO(n172), .S(n173) );
  ADDFXL U121 ( .A(b[3]), .B(b[6]), .CI(b[4]), .CO(n176), .S(n177) );
  ADDFXL U122 ( .A(b[2]), .B(b[5]), .CI(b[3]), .CO(n178), .S(n179) );
  ADDFXL U129 ( .A(b[11]), .B(b[14]), .CI(b[12]), .CO(n160), .S(n161) );
  ADDFXL U130 ( .A(b[14]), .B(b[17]), .CI(b[15]), .CO(n154), .S(n155) );
  ADDFXL U131 ( .A(b[18]), .B(b[21]), .CI(b[19]), .CO(n146), .S(n147) );
  ADDFXL U132 ( .A(b[10]), .B(b[13]), .CI(b[11]), .CO(n162), .S(n163) );
  ADDFXL U133 ( .A(b[9]), .B(b[12]), .CI(b[10]), .CO(n164), .S(n165) );
  ADDFXL U134 ( .A(b[8]), .B(b[11]), .CI(b[9]), .CO(n166), .S(n167) );
  ADDFXL U135 ( .A(b[6]), .B(b[9]), .CI(b[7]), .CO(n170), .S(n171) );
  ADDFXL U136 ( .A(b[7]), .B(b[10]), .CI(b[8]), .CO(n168), .S(n169) );
  ADDFXL U137 ( .A(b[4]), .B(b[7]), .CI(b[5]), .CO(n174), .S(n175) );
  ADDFXL U138 ( .A(b[22]), .B(b[25]), .CI(b[23]), .CO(n138), .S(n139) );
  ADDFXL U139 ( .A(b[26]), .B(b[29]), .CI(b[27]), .CO(n130), .S(n131) );
  ADDFXL U140 ( .A(b[30]), .B(b[33]), .CI(b[31]), .CO(n122), .S(n123) );
  ADDFXL U141 ( .A(b[33]), .B(b[36]), .CI(b[34]), .CO(n116), .S(n117) );
  ADDFXL U142 ( .A(b[36]), .B(b[39]), .CI(b[37]), .CO(n110), .S(n111) );
  ADDFXL U143 ( .A(b[39]), .B(b[42]), .CI(b[40]), .CO(n104), .S(n105) );
  ADDFXL U144 ( .A(b[42]), .B(b[45]), .CI(b[43]), .CO(n98), .S(n99) );
  ADDFXL U145 ( .A(b[47]), .B(b[50]), .CI(b[48]), .CO(n88), .S(n89) );
  ADDFXL U146 ( .A(b[48]), .B(b[51]), .CI(b[49]), .CO(n86), .S(n87) );
  ADDFXL U147 ( .A(b[51]), .B(b[54]), .CI(b[52]), .CO(n80), .S(n81) );
  ADDFXL U148 ( .A(n155), .B(n156), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U149 ( .A(n151), .B(n152), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U150 ( .A(n147), .B(n148), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U151 ( .A(\b[1] ), .B(b[4]), .CI(b[2]), .CO(n180), .S(n181) );
  ADDHXL U152 ( .A(b[3]), .B(\b[1] ), .CO(n182), .S(n183) );
  ADDFXL U153 ( .A(b[25]), .B(b[28]), .CI(b[26]), .CO(n132), .S(n133) );
  ADDFXL U154 ( .A(b[54]), .B(b[57]), .CI(b[55]), .CO(n74), .S(n75) );
  ADDFXL U155 ( .A(b[17]), .B(b[20]), .CI(b[18]), .CO(n148), .S(n149) );
  ADDFXL U156 ( .A(b[57]), .B(b[60]), .CI(b[58]), .CO(n68), .S(n69) );
  ADDFXL U157 ( .A(n157), .B(n158), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U158 ( .A(n177), .B(n178), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U159 ( .A(n173), .B(n174), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U160 ( .A(n169), .B(n170), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U161 ( .A(n165), .B(n166), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U162 ( .A(n161), .B(n162), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U163 ( .A(n143), .B(n144), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U164 ( .A(n139), .B(n140), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U165 ( .A(n135), .B(n136), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U166 ( .A(n131), .B(n132), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U167 ( .A(n127), .B(n128), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U168 ( .A(n123), .B(n124), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U169 ( .A(n119), .B(n120), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U170 ( .A(n115), .B(n116), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U171 ( .A(n111), .B(n112), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U172 ( .A(n107), .B(n108), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U173 ( .A(n103), .B(n104), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U174 ( .A(n99), .B(n100), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U175 ( .A(n95), .B(n96), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U176 ( .A(n91), .B(n92), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U177 ( .A(n87), .B(n88), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U178 ( .A(n83), .B(n84), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U179 ( .A(n81), .B(n82), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U180 ( .A(n79), .B(n80), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U181 ( .A(n77), .B(n78), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U182 ( .A(n75), .B(n76), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U183 ( .A(n71), .B(n72), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U184 ( .A(n67), .B(n68), .CI(n4), .CO(n3), .S(product[61]) );
  XOR2X1 U185 ( .A(n323), .B(b[63]), .Y(n321) );
  XNOR2X1 U186 ( .A(n64), .B(n2), .Y(n323) );
  ADDFXL U187 ( .A(n181), .B(n182), .CI(n61), .CO(n60), .S(product[4]) );
  ADDFXL U188 ( .A(n153), .B(n154), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U189 ( .A(n149), .B(n150), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U190 ( .A(n145), .B(n146), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U191 ( .A(n141), .B(n142), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U192 ( .A(n137), .B(n138), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U193 ( .A(n133), .B(n134), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U194 ( .A(n129), .B(n130), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U195 ( .A(n125), .B(n126), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U196 ( .A(n73), .B(n74), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U197 ( .A(n69), .B(n70), .CI(n5), .CO(n4), .S(product[60]) );
  XNOR2XL U198 ( .A(b[61]), .B(b[60]), .Y(n322) );
  XOR2X1 U199 ( .A(n321), .B(n322), .Y(product[63]) );
endmodule


module GSIM_DW_mult_tc_15 ( a, b, product );
  input [4:0] a;
  input [63:0] b;
  output [68:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, \b[0] , \b[1] , n321, n322, n323;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[1] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U4 ( .A(n67), .B(n68), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U5 ( .A(n69), .B(n70), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U12 ( .A(n83), .B(n84), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U14 ( .A(n87), .B(n88), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U16 ( .A(n91), .B(n92), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U18 ( .A(n95), .B(n96), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U20 ( .A(n99), .B(n100), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U22 ( .A(n103), .B(n104), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U24 ( .A(n107), .B(n108), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U26 ( .A(n111), .B(n112), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U28 ( .A(n115), .B(n116), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U49 ( .A(n157), .B(n158), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U52 ( .A(n163), .B(n164), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U54 ( .A(n167), .B(n168), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U56 ( .A(n171), .B(n172), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U58 ( .A(n175), .B(n176), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U61 ( .A(n181), .B(n182), .CI(n61), .CO(n60), .S(product[4]) );
  ADDFXL U66 ( .A(b[58]), .B(b[61]), .CI(b[59]), .CO(n66), .S(n67) );
  ADDFXL U67 ( .A(b[57]), .B(b[60]), .CI(b[58]), .CO(n68), .S(n69) );
  ADDFXL U69 ( .A(b[55]), .B(b[58]), .CI(b[56]), .CO(n72), .S(n73) );
  ADDFXL U70 ( .A(b[54]), .B(b[57]), .CI(b[55]), .CO(n74), .S(n75) );
  ADDFXL U72 ( .A(b[52]), .B(b[55]), .CI(b[53]), .CO(n78), .S(n79) );
  ADDFXL U73 ( .A(b[51]), .B(b[54]), .CI(b[52]), .CO(n80), .S(n81) );
  ADDFXL U75 ( .A(b[49]), .B(b[52]), .CI(b[50]), .CO(n84), .S(n85) );
  ADDFXL U76 ( .A(b[48]), .B(b[51]), .CI(b[49]), .CO(n86), .S(n87) );
  ADDFXL U78 ( .A(b[46]), .B(b[49]), .CI(b[47]), .CO(n90), .S(n91) );
  ADDFXL U79 ( .A(b[45]), .B(b[48]), .CI(b[46]), .CO(n92), .S(n93) );
  ADDFXL U81 ( .A(b[43]), .B(b[46]), .CI(b[44]), .CO(n96), .S(n97) );
  ADDFXL U82 ( .A(b[42]), .B(b[45]), .CI(b[43]), .CO(n98), .S(n99) );
  ADDFXL U85 ( .A(b[39]), .B(b[42]), .CI(b[40]), .CO(n104), .S(n105) );
  ADDFXL U86 ( .A(b[38]), .B(b[41]), .CI(b[39]), .CO(n106), .S(n107) );
  ADDFXL U88 ( .A(b[36]), .B(b[39]), .CI(b[37]), .CO(n110), .S(n111) );
  ADDFXL U89 ( .A(b[35]), .B(b[38]), .CI(b[36]), .CO(n112), .S(n113) );
  ADDFXL U91 ( .A(b[33]), .B(b[36]), .CI(b[34]), .CO(n116), .S(n117) );
  ADDFXL U92 ( .A(b[32]), .B(b[35]), .CI(b[33]), .CO(n118), .S(n119) );
  ADDFXL U94 ( .A(b[30]), .B(b[33]), .CI(b[31]), .CO(n122), .S(n123) );
  ADDFXL U95 ( .A(b[29]), .B(b[32]), .CI(b[30]), .CO(n124), .S(n125) );
  ADDFXL U97 ( .A(b[27]), .B(b[30]), .CI(b[28]), .CO(n128), .S(n129) );
  ADDFXL U98 ( .A(b[26]), .B(b[29]), .CI(b[27]), .CO(n130), .S(n131) );
  ADDFXL U101 ( .A(b[23]), .B(b[26]), .CI(b[24]), .CO(n136), .S(n137) );
  ADDFXL U102 ( .A(b[22]), .B(b[25]), .CI(b[23]), .CO(n138), .S(n139) );
  ADDFXL U104 ( .A(b[20]), .B(b[23]), .CI(b[21]), .CO(n142), .S(n143) );
  ADDFXL U105 ( .A(b[19]), .B(b[22]), .CI(b[20]), .CO(n144), .S(n145) );
  ADDFXL U108 ( .A(b[16]), .B(b[19]), .CI(b[17]), .CO(n150), .S(n151) );
  ADDFXL U111 ( .A(b[13]), .B(b[16]), .CI(b[14]), .CO(n156), .S(n157) );
  ADDFXL U114 ( .A(b[10]), .B(b[13]), .CI(b[11]), .CO(n162), .S(n163) );
  ADDFXL U117 ( .A(b[7]), .B(b[10]), .CI(b[8]), .CO(n168), .S(n169) );
  ADDFXL U119 ( .A(b[5]), .B(b[8]), .CI(b[6]), .CO(n172), .S(n173) );
  ADDFXL U120 ( .A(b[4]), .B(b[7]), .CI(b[5]), .CO(n174), .S(n175) );
  ADDFXL U129 ( .A(b[6]), .B(b[9]), .CI(b[7]), .CO(n170), .S(n171) );
  ADDFXL U130 ( .A(b[8]), .B(b[11]), .CI(b[9]), .CO(n166), .S(n167) );
  ADDFXL U131 ( .A(b[11]), .B(b[14]), .CI(b[12]), .CO(n160), .S(n161) );
  ADDFXL U132 ( .A(b[14]), .B(b[17]), .CI(b[15]), .CO(n154), .S(n155) );
  ADDFXL U133 ( .A(b[17]), .B(b[20]), .CI(b[18]), .CO(n148), .S(n149) );
  ADDFXL U134 ( .A(b[2]), .B(b[5]), .CI(b[3]), .CO(n178), .S(n179) );
  ADDFHX2 U135 ( .A(\b[1] ), .B(b[4]), .CI(b[2]), .CO(n180), .S(n181) );
  ADDHXL U136 ( .A(b[3]), .B(\b[1] ), .CO(n182), .S(n183) );
  ADDFX2 U137 ( .A(n62), .B(\b[0] ), .CI(n183), .CO(n61), .S(product[3]) );
  ADDFXL U138 ( .A(b[9]), .B(b[12]), .CI(b[10]), .CO(n164), .S(n165) );
  ADDFXL U139 ( .A(b[12]), .B(b[15]), .CI(b[13]), .CO(n158), .S(n159) );
  ADDFXL U140 ( .A(b[15]), .B(b[18]), .CI(b[16]), .CO(n152), .S(n153) );
  ADDFXL U141 ( .A(b[18]), .B(b[21]), .CI(b[19]), .CO(n146), .S(n147) );
  ADDFXL U142 ( .A(b[21]), .B(b[24]), .CI(b[22]), .CO(n140), .S(n141) );
  ADDFXL U143 ( .A(b[25]), .B(b[28]), .CI(b[26]), .CO(n132), .S(n133) );
  ADDFXL U144 ( .A(b[31]), .B(b[34]), .CI(b[32]), .CO(n120), .S(n121) );
  ADDFXL U145 ( .A(b[34]), .B(b[37]), .CI(b[35]), .CO(n114), .S(n115) );
  ADDFXL U146 ( .A(b[37]), .B(b[40]), .CI(b[38]), .CO(n108), .S(n109) );
  ADDFXL U147 ( .A(b[41]), .B(b[44]), .CI(b[42]), .CO(n100), .S(n101) );
  ADDFXL U148 ( .A(b[44]), .B(b[47]), .CI(b[45]), .CO(n94), .S(n95) );
  ADDFXL U149 ( .A(b[47]), .B(b[50]), .CI(b[48]), .CO(n88), .S(n89) );
  ADDFXL U150 ( .A(b[50]), .B(b[53]), .CI(b[51]), .CO(n82), .S(n83) );
  ADDFXL U151 ( .A(b[24]), .B(b[27]), .CI(b[25]), .CO(n134), .S(n135) );
  ADDFXL U152 ( .A(b[59]), .B(b[62]), .CI(b[60]), .CO(n64), .S(n65) );
  ADDFXL U153 ( .A(b[28]), .B(b[31]), .CI(b[29]), .CO(n126), .S(n127) );
  ADDFXL U154 ( .A(b[40]), .B(b[43]), .CI(b[41]), .CO(n102), .S(n103) );
  ADDFXL U155 ( .A(b[56]), .B(b[59]), .CI(b[57]), .CO(n70), .S(n71) );
  ADDFXL U156 ( .A(b[53]), .B(b[56]), .CI(b[54]), .CO(n76), .S(n77) );
  CMPR32X2 U157 ( .A(b[3]), .B(b[6]), .C(b[4]), .CO(n176), .S(n177) );
  ADDHX2 U158 ( .A(\b[0] ), .B(b[2]), .CO(n62), .S(product[2]) );
  ADDFXL U159 ( .A(n179), .B(n180), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U160 ( .A(n177), .B(n178), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U161 ( .A(n169), .B(n170), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U162 ( .A(n165), .B(n166), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U163 ( .A(n173), .B(n174), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U164 ( .A(n159), .B(n160), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U165 ( .A(n155), .B(n156), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U166 ( .A(n161), .B(n162), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U167 ( .A(n147), .B(n148), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U168 ( .A(n149), .B(n150), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U169 ( .A(n151), .B(n152), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U170 ( .A(n153), .B(n154), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U171 ( .A(n141), .B(n142), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U172 ( .A(n143), .B(n144), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U173 ( .A(n145), .B(n146), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U174 ( .A(n135), .B(n136), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U175 ( .A(n137), .B(n138), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U176 ( .A(n139), .B(n140), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U177 ( .A(n127), .B(n128), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U178 ( .A(n129), .B(n130), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U179 ( .A(n131), .B(n132), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U180 ( .A(n133), .B(n134), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U181 ( .A(n121), .B(n122), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U182 ( .A(n123), .B(n124), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U183 ( .A(n125), .B(n126), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U184 ( .A(n117), .B(n118), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U185 ( .A(n113), .B(n114), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U186 ( .A(n109), .B(n110), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U187 ( .A(n105), .B(n106), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U188 ( .A(n101), .B(n102), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U189 ( .A(n97), .B(n98), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U190 ( .A(n93), .B(n94), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U191 ( .A(n89), .B(n90), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U192 ( .A(n85), .B(n86), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U193 ( .A(n79), .B(n80), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U194 ( .A(n77), .B(n78), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U195 ( .A(n65), .B(n66), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U196 ( .A(n73), .B(n74), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U197 ( .A(n119), .B(n120), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U198 ( .A(n81), .B(n82), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U199 ( .A(n75), .B(n76), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U200 ( .A(n71), .B(n72), .CI(n6), .CO(n5), .S(product[59]) );
  XNOR2XL U201 ( .A(b[61]), .B(b[60]), .Y(n322) );
  XOR2X1 U202 ( .A(n321), .B(n322), .Y(product[63]) );
  XOR2X1 U203 ( .A(n323), .B(b[63]), .Y(n321) );
  XNOR2X1 U204 ( .A(n64), .B(n2), .Y(n323) );
endmodule


module GSIM_DW01_add_494 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;
  assign SUM[0] = B[0];

  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  XOR3X2 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2XL U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module GSIM_DW01_add_493 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module GSIM_DW01_add_492 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFHX2 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module GSIM_DW_mult_tc_14 ( a, b, product );
  input [3:0] a;
  input [63:0] b;
  output [67:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, \b[0] , \b[1] , n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318;
  assign product[1] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[2] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U4 ( .A(b[60]), .B(n316), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U5 ( .A(b[59]), .B(n315), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U6 ( .A(b[58]), .B(n314), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U7 ( .A(b[57]), .B(n313), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U8 ( .A(b[56]), .B(n312), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U9 ( .A(b[55]), .B(n311), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U10 ( .A(b[54]), .B(n310), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U11 ( .A(b[53]), .B(n309), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U14 ( .A(b[50]), .B(n306), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U15 ( .A(b[49]), .B(n305), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U16 ( .A(b[48]), .B(n304), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U17 ( .A(b[47]), .B(n303), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U18 ( .A(b[46]), .B(n302), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U19 ( .A(b[45]), .B(n301), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U20 ( .A(b[44]), .B(n300), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U21 ( .A(b[43]), .B(n299), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U24 ( .A(b[40]), .B(n296), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U25 ( .A(b[39]), .B(n295), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U26 ( .A(b[38]), .B(n294), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U27 ( .A(b[37]), .B(n293), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U28 ( .A(b[36]), .B(n292), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U29 ( .A(b[35]), .B(n291), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U30 ( .A(b[34]), .B(n290), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U31 ( .A(b[33]), .B(n289), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U34 ( .A(b[30]), .B(n286), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U35 ( .A(b[29]), .B(n285), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U36 ( .A(b[28]), .B(n284), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U37 ( .A(b[27]), .B(n283), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U38 ( .A(b[26]), .B(n282), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U39 ( .A(b[25]), .B(n281), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U40 ( .A(b[24]), .B(n280), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U41 ( .A(b[23]), .B(n279), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U44 ( .A(b[20]), .B(n276), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U45 ( .A(b[19]), .B(n275), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U46 ( .A(b[18]), .B(n274), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U47 ( .A(b[17]), .B(n273), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U48 ( .A(b[16]), .B(n272), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U49 ( .A(b[15]), .B(n271), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U50 ( .A(b[14]), .B(n270), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U51 ( .A(b[13]), .B(n269), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U54 ( .A(b[10]), .B(n266), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U55 ( .A(b[9]), .B(n265), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U56 ( .A(b[8]), .B(n264), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U57 ( .A(b[7]), .B(n263), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U58 ( .A(b[6]), .B(n262), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U59 ( .A(b[5]), .B(n261), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U131 ( .A(b[31]), .B(n287), .CI(n33), .CO(n32), .S(product[32]) );
  CLKINVX1 U132 ( .A(b[3]), .Y(n261) );
  ADDFXL U133 ( .A(b[3]), .B(n259), .CI(n61), .CO(n60), .S(product[4]) );
  ADDFXL U134 ( .A(b[22]), .B(n278), .CI(n42), .CO(n41), .S(product[23]) );
  XOR2XL U135 ( .A(b[2]), .B(\b[0] ), .Y(product[3]) );
  ADDFXL U136 ( .A(b[41]), .B(n297), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U137 ( .A(b[61]), .B(n317), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U138 ( .A(b[52]), .B(n308), .CI(n12), .CO(n11), .S(product[53]) );
  INVX1 U139 ( .A(\b[1] ), .Y(n259) );
  INVXL U140 ( .A(b[16]), .Y(n274) );
  INVXL U141 ( .A(b[28]), .Y(n286) );
  INVXL U142 ( .A(b[36]), .Y(n294) );
  INVXL U143 ( .A(b[48]), .Y(n306) );
  INVXL U144 ( .A(b[8]), .Y(n266) );
  INVXL U145 ( .A(b[18]), .Y(n276) );
  INVXL U146 ( .A(b[38]), .Y(n296) );
  INVXL U147 ( .A(b[12]), .Y(n270) );
  INVXL U148 ( .A(b[22]), .Y(n280) );
  INVXL U149 ( .A(b[32]), .Y(n290) );
  INVXL U150 ( .A(b[42]), .Y(n300) );
  INVXL U151 ( .A(b[4]), .Y(n262) );
  INVXL U152 ( .A(b[11]), .Y(n269) );
  INVXL U153 ( .A(b[21]), .Y(n279) );
  INVXL U154 ( .A(b[31]), .Y(n289) );
  INVXL U155 ( .A(b[41]), .Y(n299) );
  INVXL U156 ( .A(b[14]), .Y(n272) );
  INVXL U157 ( .A(b[24]), .Y(n282) );
  INVXL U158 ( .A(b[34]), .Y(n292) );
  INVXL U159 ( .A(b[44]), .Y(n302) );
  INVXL U160 ( .A(b[5]), .Y(n263) );
  INVXL U161 ( .A(b[6]), .Y(n264) );
  INVXL U162 ( .A(b[7]), .Y(n265) );
  INVXL U163 ( .A(b[13]), .Y(n271) );
  INVXL U164 ( .A(b[15]), .Y(n273) );
  INVXL U165 ( .A(b[17]), .Y(n275) );
  INVXL U166 ( .A(b[23]), .Y(n281) );
  INVXL U167 ( .A(b[25]), .Y(n283) );
  INVXL U168 ( .A(b[26]), .Y(n284) );
  INVXL U169 ( .A(b[27]), .Y(n285) );
  INVXL U170 ( .A(b[33]), .Y(n291) );
  INVXL U171 ( .A(b[35]), .Y(n293) );
  INVXL U172 ( .A(b[37]), .Y(n295) );
  INVXL U173 ( .A(b[43]), .Y(n301) );
  INVXL U174 ( .A(b[45]), .Y(n303) );
  INVXL U175 ( .A(b[46]), .Y(n304) );
  INVXL U176 ( .A(b[47]), .Y(n305) );
  INVXL U177 ( .A(b[2]), .Y(n260) );
  ADDFXL U178 ( .A(b[11]), .B(n267), .CI(n53), .CO(n52), .S(product[12]) );
  INVXL U179 ( .A(b[9]), .Y(n267) );
  ADDFXL U180 ( .A(b[21]), .B(n277), .CI(n43), .CO(n42), .S(product[22]) );
  INVXL U181 ( .A(b[19]), .Y(n277) );
  INVXL U182 ( .A(b[29]), .Y(n287) );
  INVXL U183 ( .A(b[39]), .Y(n297) );
  ADDFXL U184 ( .A(b[4]), .B(n260), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U185 ( .A(b[12]), .B(n268), .CI(n52), .CO(n51), .S(product[13]) );
  INVXL U186 ( .A(b[10]), .Y(n268) );
  INVXL U187 ( .A(b[20]), .Y(n278) );
  ADDFXL U188 ( .A(b[32]), .B(n288), .CI(n32), .CO(n31), .S(product[33]) );
  INVXL U189 ( .A(b[30]), .Y(n288) );
  ADDFXL U190 ( .A(b[42]), .B(n298), .CI(n22), .CO(n21), .S(product[43]) );
  INVXL U191 ( .A(b[40]), .Y(n298) );
  INVXL U192 ( .A(b[58]), .Y(n316) );
  INVXL U193 ( .A(b[52]), .Y(n310) );
  INVXL U194 ( .A(b[51]), .Y(n309) );
  INVXL U195 ( .A(b[54]), .Y(n312) );
  INVXL U196 ( .A(b[53]), .Y(n311) );
  INVXL U197 ( .A(b[55]), .Y(n313) );
  INVXL U198 ( .A(b[56]), .Y(n314) );
  INVXL U199 ( .A(b[57]), .Y(n315) );
  ADDFXL U200 ( .A(b[51]), .B(n307), .CI(n13), .CO(n12), .S(product[52]) );
  INVXL U201 ( .A(b[49]), .Y(n307) );
  INVXL U202 ( .A(b[59]), .Y(n317) );
  INVXL U203 ( .A(b[50]), .Y(n308) );
  XOR2X1 U204 ( .A(n318), .B(b[60]), .Y(product[63]) );
  XNOR2X1 U205 ( .A(n2), .B(b[62]), .Y(n318) );
  NAND2X1 U206 ( .A(\b[0] ), .B(n260), .Y(n61) );
endmodule


module GSIM_DW01_add_491 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;
  assign SUM[15] = B[15];
  assign SUM[14] = B[14];
  assign SUM[13] = B[13];
  assign SUM[12] = B[12];
  assign SUM[11] = B[11];
  assign SUM[10] = B[10];
  assign SUM[9] = B[9];
  assign SUM[8] = B[8];
  assign SUM[7] = B[7];
  assign SUM[6] = B[6];
  assign SUM[5] = B[5];
  assign SUM[4] = B[4];
  assign SUM[3] = B[3];
  assign SUM[2] = B[2];
  assign SUM[1] = B[1];

  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(n1), .CO(carry[18]), .S(SUM[17]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  XOR3X2 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  AND2X2 U1 ( .A(B[16]), .B(A[16]), .Y(n1) );
  XOR2XL U2 ( .A(B[16]), .B(A[16]), .Y(SUM[16]) );
endmodule


module GSIM_DW_mult_tc_13 ( a, b, product );
  input [4:0] a;
  input [63:0] b;
  output [68:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, \b[0] , \b[1] , n321, n322, n323;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[1] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U4 ( .A(n67), .B(n68), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U15 ( .A(n89), .B(n90), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U17 ( .A(n93), .B(n94), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U19 ( .A(n97), .B(n98), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U25 ( .A(n109), .B(n110), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U27 ( .A(n113), .B(n114), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U29 ( .A(n117), .B(n118), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U49 ( .A(n157), .B(n158), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U55 ( .A(n169), .B(n170), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U57 ( .A(n173), .B(n174), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U62 ( .A(n62), .B(\b[0] ), .CI(n183), .CO(n61), .S(product[3]) );
  ADDFXL U65 ( .A(b[59]), .B(b[62]), .CI(b[60]), .CO(n64), .S(n65) );
  ADDFXL U66 ( .A(b[58]), .B(b[61]), .CI(b[59]), .CO(n66), .S(n67) );
  ADDFXL U68 ( .A(b[56]), .B(b[59]), .CI(b[57]), .CO(n70), .S(n71) );
  ADDFXL U69 ( .A(b[55]), .B(b[58]), .CI(b[56]), .CO(n72), .S(n73) );
  ADDFXL U71 ( .A(b[53]), .B(b[56]), .CI(b[54]), .CO(n76), .S(n77) );
  ADDFXL U72 ( .A(b[52]), .B(b[55]), .CI(b[53]), .CO(n78), .S(n79) );
  ADDFXL U74 ( .A(b[50]), .B(b[53]), .CI(b[51]), .CO(n82), .S(n83) );
  ADDFXL U75 ( .A(b[49]), .B(b[52]), .CI(b[50]), .CO(n84), .S(n85) );
  ADDFXL U78 ( .A(b[46]), .B(b[49]), .CI(b[47]), .CO(n90), .S(n91) );
  ADDFXL U79 ( .A(b[45]), .B(b[48]), .CI(b[46]), .CO(n92), .S(n93) );
  ADDFXL U80 ( .A(b[44]), .B(b[47]), .CI(b[45]), .CO(n94), .S(n95) );
  ADDFXL U81 ( .A(b[43]), .B(b[46]), .CI(b[44]), .CO(n96), .S(n97) );
  ADDFXL U83 ( .A(b[41]), .B(b[44]), .CI(b[42]), .CO(n100), .S(n101) );
  ADDFXL U84 ( .A(b[40]), .B(b[43]), .CI(b[41]), .CO(n102), .S(n103) );
  ADDFXL U86 ( .A(b[38]), .B(b[41]), .CI(b[39]), .CO(n106), .S(n107) );
  ADDFXL U87 ( .A(b[37]), .B(b[40]), .CI(b[38]), .CO(n108), .S(n109) );
  ADDFXL U89 ( .A(b[35]), .B(b[38]), .CI(b[36]), .CO(n112), .S(n113) );
  ADDFXL U90 ( .A(b[34]), .B(b[37]), .CI(b[35]), .CO(n114), .S(n115) );
  ADDFXL U92 ( .A(b[32]), .B(b[35]), .CI(b[33]), .CO(n118), .S(n119) );
  ADDFXL U93 ( .A(b[31]), .B(b[34]), .CI(b[32]), .CO(n120), .S(n121) );
  ADDFXL U95 ( .A(b[29]), .B(b[32]), .CI(b[30]), .CO(n124), .S(n125) );
  ADDFXL U96 ( .A(b[28]), .B(b[31]), .CI(b[29]), .CO(n126), .S(n127) );
  ADDFXL U97 ( .A(b[27]), .B(b[30]), .CI(b[28]), .CO(n128), .S(n129) );
  ADDFXL U100 ( .A(b[24]), .B(b[27]), .CI(b[25]), .CO(n134), .S(n135) );
  ADDFXL U101 ( .A(b[23]), .B(b[26]), .CI(b[24]), .CO(n136), .S(n137) );
  ADDFXL U103 ( .A(b[21]), .B(b[24]), .CI(b[22]), .CO(n140), .S(n141) );
  ADDFXL U104 ( .A(b[20]), .B(b[23]), .CI(b[21]), .CO(n142), .S(n143) );
  ADDFXL U105 ( .A(b[19]), .B(b[22]), .CI(b[20]), .CO(n144), .S(n145) );
  ADDFXL U108 ( .A(b[16]), .B(b[19]), .CI(b[17]), .CO(n150), .S(n151) );
  ADDFXL U109 ( .A(b[15]), .B(b[18]), .CI(b[16]), .CO(n152), .S(n153) );
  ADDFXL U111 ( .A(b[13]), .B(b[16]), .CI(b[14]), .CO(n156), .S(n157) );
  ADDFXL U112 ( .A(b[12]), .B(b[15]), .CI(b[13]), .CO(n158), .S(n159) );
  ADDFXL U114 ( .A(b[10]), .B(b[13]), .CI(b[11]), .CO(n162), .S(n163) );
  ADDFXL U119 ( .A(b[5]), .B(b[8]), .CI(b[6]), .CO(n172), .S(n173) );
  ADDFXL U121 ( .A(b[3]), .B(b[6]), .CI(b[4]), .CO(n176), .S(n177) );
  ADDFXL U129 ( .A(b[9]), .B(b[12]), .CI(b[10]), .CO(n164), .S(n165) );
  ADDFXL U130 ( .A(b[8]), .B(b[11]), .CI(b[9]), .CO(n166), .S(n167) );
  ADDFXL U131 ( .A(b[6]), .B(b[9]), .CI(b[7]), .CO(n170), .S(n171) );
  ADDFXL U132 ( .A(b[7]), .B(b[10]), .CI(b[8]), .CO(n168), .S(n169) );
  ADDFXL U133 ( .A(b[4]), .B(b[7]), .CI(b[5]), .CO(n174), .S(n175) );
  ADDHXL U134 ( .A(b[3]), .B(\b[1] ), .CO(n182), .S(n183) );
  ADDFXL U135 ( .A(n181), .B(n182), .CI(n61), .CO(n60), .S(product[4]) );
  ADDFXL U136 ( .A(b[14]), .B(b[17]), .CI(b[15]), .CO(n154), .S(n155) );
  ADDFXL U137 ( .A(b[18]), .B(b[21]), .CI(b[19]), .CO(n146), .S(n147) );
  ADDFXL U138 ( .A(b[22]), .B(b[25]), .CI(b[23]), .CO(n138), .S(n139) );
  ADDFXL U139 ( .A(b[26]), .B(b[29]), .CI(b[27]), .CO(n130), .S(n131) );
  ADDFXL U140 ( .A(b[30]), .B(b[33]), .CI(b[31]), .CO(n122), .S(n123) );
  ADDFXL U141 ( .A(b[33]), .B(b[36]), .CI(b[34]), .CO(n116), .S(n117) );
  ADDFXL U142 ( .A(b[36]), .B(b[39]), .CI(b[37]), .CO(n110), .S(n111) );
  ADDFXL U143 ( .A(b[39]), .B(b[42]), .CI(b[40]), .CO(n104), .S(n105) );
  ADDFXL U144 ( .A(b[42]), .B(b[45]), .CI(b[43]), .CO(n98), .S(n99) );
  ADDFXL U145 ( .A(b[48]), .B(b[51]), .CI(b[49]), .CO(n86), .S(n87) );
  ADDFXL U146 ( .A(b[51]), .B(b[54]), .CI(b[52]), .CO(n80), .S(n81) );
  ADDFXL U147 ( .A(b[47]), .B(b[50]), .CI(b[48]), .CO(n88), .S(n89) );
  ADDFXL U148 ( .A(b[25]), .B(b[28]), .CI(b[26]), .CO(n132), .S(n133) );
  ADDFXL U149 ( .A(b[54]), .B(b[57]), .CI(b[55]), .CO(n74), .S(n75) );
  ADDFXL U150 ( .A(b[17]), .B(b[20]), .CI(b[18]), .CO(n148), .S(n149) );
  ADDFXL U151 ( .A(b[11]), .B(b[14]), .CI(b[12]), .CO(n160), .S(n161) );
  ADDFXL U152 ( .A(b[57]), .B(b[60]), .CI(b[58]), .CO(n68), .S(n69) );
  ADDFXL U153 ( .A(b[2]), .B(b[5]), .CI(b[3]), .CO(n178), .S(n179) );
  ADDFXL U154 ( .A(n171), .B(n172), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U155 ( .A(n167), .B(n168), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U156 ( .A(n159), .B(n160), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U157 ( .A(n163), .B(n164), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U158 ( .A(n155), .B(n156), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U159 ( .A(n153), .B(n154), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U160 ( .A(n143), .B(n144), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U161 ( .A(n149), .B(n150), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U162 ( .A(n141), .B(n142), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U163 ( .A(n147), .B(n148), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U164 ( .A(n135), .B(n136), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U165 ( .A(n137), .B(n138), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U166 ( .A(n139), .B(n140), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U167 ( .A(n127), .B(n128), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U168 ( .A(n131), .B(n132), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U169 ( .A(n123), .B(n124), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U170 ( .A(n119), .B(n120), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U171 ( .A(n115), .B(n116), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U172 ( .A(n111), .B(n112), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U173 ( .A(n107), .B(n108), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U174 ( .A(n103), .B(n104), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U175 ( .A(n99), .B(n100), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U176 ( .A(n95), .B(n96), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U177 ( .A(n91), .B(n92), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U178 ( .A(n83), .B(n84), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U179 ( .A(n77), .B(n78), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U180 ( .A(n73), .B(n74), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U181 ( .A(n87), .B(n88), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U182 ( .A(n69), .B(n70), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U183 ( .A(n65), .B(n66), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U184 ( .A(\b[1] ), .B(b[4]), .CI(b[2]), .CO(n180), .S(n181) );
  XOR2X1 U185 ( .A(n321), .B(n322), .Y(product[63]) );
  ADDHX1 U186 ( .A(\b[0] ), .B(b[2]), .CO(n62), .S(product[2]) );
  ADDFX1 U187 ( .A(n179), .B(n180), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U188 ( .A(n175), .B(n176), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U189 ( .A(n151), .B(n152), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U190 ( .A(n145), .B(n146), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U191 ( .A(n133), .B(n134), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U192 ( .A(n129), .B(n130), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U193 ( .A(n125), .B(n126), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U194 ( .A(n121), .B(n122), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U195 ( .A(n79), .B(n80), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U196 ( .A(n71), .B(n72), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U197 ( .A(n75), .B(n76), .CI(n8), .CO(n7), .S(product[57]) );
  XNOR2XL U198 ( .A(b[61]), .B(b[60]), .Y(n322) );
  ADDFXL U199 ( .A(n165), .B(n166), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U200 ( .A(n177), .B(n178), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U201 ( .A(n161), .B(n162), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U202 ( .A(n105), .B(n106), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U203 ( .A(n85), .B(n86), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U204 ( .A(n101), .B(n102), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U205 ( .A(n81), .B(n82), .CI(n11), .CO(n10), .S(product[54]) );
  XOR2X1 U206 ( .A(n323), .B(b[63]), .Y(n321) );
  XNOR2X1 U207 ( .A(n64), .B(n2), .Y(n323) );
endmodule


module GSIM_DW01_add_490 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;
  assign SUM[0] = B[0];

  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR3X2 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2XL U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module GSIM_DW01_add_489 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;

  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XL U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module GSIM_DW_mult_tc_5 ( a, b, product );
  input [4:0] a;
  input [63:0] b;
  output [68:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, \b[0] , \b[1] , n321, n322, n323;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[1] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U4 ( .A(n67), .B(n68), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U11 ( .A(n81), .B(n82), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U13 ( .A(n85), .B(n86), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U15 ( .A(n89), .B(n90), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U17 ( .A(n93), .B(n94), .CI(n17), .CO(n16), .S(product[48]) );
  ADDFXL U21 ( .A(n101), .B(n102), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U23 ( .A(n105), .B(n106), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U25 ( .A(n109), .B(n110), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U27 ( .A(n113), .B(n114), .CI(n27), .CO(n26), .S(product[38]) );
  ADDFXL U31 ( .A(n121), .B(n122), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U51 ( .A(n161), .B(n162), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U53 ( .A(n165), .B(n166), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U55 ( .A(n169), .B(n170), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U57 ( .A(n173), .B(n174), .CI(n57), .CO(n56), .S(product[8]) );
  ADDFXL U61 ( .A(n181), .B(n182), .CI(n61), .CO(n60), .S(product[4]) );
  ADDFXL U66 ( .A(b[58]), .B(b[61]), .CI(b[59]), .CO(n66), .S(n67) );
  ADDFXL U67 ( .A(b[57]), .B(b[60]), .CI(b[58]), .CO(n68), .S(n69) );
  ADDFXL U69 ( .A(b[55]), .B(b[58]), .CI(b[56]), .CO(n72), .S(n73) );
  ADDFXL U70 ( .A(b[54]), .B(b[57]), .CI(b[55]), .CO(n74), .S(n75) );
  ADDFXL U72 ( .A(b[52]), .B(b[55]), .CI(b[53]), .CO(n78), .S(n79) );
  ADDFXL U73 ( .A(b[51]), .B(b[54]), .CI(b[52]), .CO(n80), .S(n81) );
  ADDFXL U75 ( .A(b[49]), .B(b[52]), .CI(b[50]), .CO(n84), .S(n85) );
  ADDFXL U76 ( .A(b[48]), .B(b[51]), .CI(b[49]), .CO(n86), .S(n87) );
  ADDFXL U78 ( .A(b[46]), .B(b[49]), .CI(b[47]), .CO(n90), .S(n91) );
  ADDFXL U79 ( .A(b[45]), .B(b[48]), .CI(b[46]), .CO(n92), .S(n93) );
  ADDFXL U81 ( .A(b[43]), .B(b[46]), .CI(b[44]), .CO(n96), .S(n97) );
  ADDFXL U82 ( .A(b[42]), .B(b[45]), .CI(b[43]), .CO(n98), .S(n99) );
  ADDFXL U85 ( .A(b[39]), .B(b[42]), .CI(b[40]), .CO(n104), .S(n105) );
  ADDFXL U86 ( .A(b[38]), .B(b[41]), .CI(b[39]), .CO(n106), .S(n107) );
  ADDFXL U88 ( .A(b[36]), .B(b[39]), .CI(b[37]), .CO(n110), .S(n111) );
  ADDFXL U89 ( .A(b[35]), .B(b[38]), .CI(b[36]), .CO(n112), .S(n113) );
  ADDFXL U91 ( .A(b[33]), .B(b[36]), .CI(b[34]), .CO(n116), .S(n117) );
  ADDFXL U92 ( .A(b[32]), .B(b[35]), .CI(b[33]), .CO(n118), .S(n119) );
  ADDFXL U94 ( .A(b[30]), .B(b[33]), .CI(b[31]), .CO(n122), .S(n123) );
  ADDFXL U95 ( .A(b[29]), .B(b[32]), .CI(b[30]), .CO(n124), .S(n125) );
  ADDFXL U97 ( .A(b[27]), .B(b[30]), .CI(b[28]), .CO(n128), .S(n129) );
  ADDFXL U98 ( .A(b[26]), .B(b[29]), .CI(b[27]), .CO(n130), .S(n131) );
  ADDFXL U101 ( .A(b[23]), .B(b[26]), .CI(b[24]), .CO(n136), .S(n137) );
  ADDFXL U102 ( .A(b[22]), .B(b[25]), .CI(b[23]), .CO(n138), .S(n139) );
  ADDFXL U104 ( .A(b[20]), .B(b[23]), .CI(b[21]), .CO(n142), .S(n143) );
  ADDFXL U105 ( .A(b[19]), .B(b[22]), .CI(b[20]), .CO(n144), .S(n145) );
  ADDFXL U108 ( .A(b[16]), .B(b[19]), .CI(b[17]), .CO(n150), .S(n151) );
  ADDFXL U110 ( .A(b[14]), .B(b[17]), .CI(b[15]), .CO(n154), .S(n155) );
  ADDFXL U111 ( .A(b[13]), .B(b[16]), .CI(b[14]), .CO(n156), .S(n157) );
  ADDFXL U114 ( .A(b[10]), .B(b[13]), .CI(b[11]), .CO(n162), .S(n163) );
  ADDFXL U117 ( .A(b[7]), .B(b[10]), .CI(b[8]), .CO(n168), .S(n169) );
  ADDFXL U119 ( .A(b[5]), .B(b[8]), .CI(b[6]), .CO(n172), .S(n173) );
  ADDFXL U120 ( .A(b[4]), .B(b[7]), .CI(b[5]), .CO(n174), .S(n175) );
  ADDFXL U121 ( .A(b[3]), .B(b[6]), .CI(b[4]), .CO(n176), .S(n177) );
  ADDFXL U129 ( .A(b[6]), .B(b[9]), .CI(b[7]), .CO(n170), .S(n171) );
  ADDFX1 U130 ( .A(\b[1] ), .B(b[4]), .CI(b[2]), .CO(n180), .S(n181) );
  ADDFXL U131 ( .A(b[8]), .B(b[11]), .CI(b[9]), .CO(n166), .S(n167) );
  ADDFXL U132 ( .A(b[11]), .B(b[14]), .CI(b[12]), .CO(n160), .S(n161) );
  ADDFXL U133 ( .A(b[17]), .B(b[20]), .CI(b[18]), .CO(n148), .S(n149) );
  ADDFXL U134 ( .A(b[2]), .B(b[5]), .CI(b[3]), .CO(n178), .S(n179) );
  ADDHXL U135 ( .A(b[3]), .B(\b[1] ), .CO(n182), .S(n183) );
  ADDFXL U136 ( .A(n62), .B(\b[0] ), .CI(n183), .CO(n61), .S(product[3]) );
  ADDFXL U137 ( .A(b[9]), .B(b[12]), .CI(b[10]), .CO(n164), .S(n165) );
  ADDFXL U138 ( .A(b[12]), .B(b[15]), .CI(b[13]), .CO(n158), .S(n159) );
  ADDFXL U139 ( .A(b[15]), .B(b[18]), .CI(b[16]), .CO(n152), .S(n153) );
  ADDFXL U140 ( .A(b[18]), .B(b[21]), .CI(b[19]), .CO(n146), .S(n147) );
  ADDFXL U141 ( .A(b[21]), .B(b[24]), .CI(b[22]), .CO(n140), .S(n141) );
  ADDFXL U142 ( .A(b[25]), .B(b[28]), .CI(b[26]), .CO(n132), .S(n133) );
  ADDFXL U143 ( .A(b[31]), .B(b[34]), .CI(b[32]), .CO(n120), .S(n121) );
  ADDFXL U144 ( .A(b[34]), .B(b[37]), .CI(b[35]), .CO(n114), .S(n115) );
  ADDFXL U145 ( .A(b[37]), .B(b[40]), .CI(b[38]), .CO(n108), .S(n109) );
  ADDFXL U146 ( .A(b[41]), .B(b[44]), .CI(b[42]), .CO(n100), .S(n101) );
  ADDFXL U147 ( .A(b[44]), .B(b[47]), .CI(b[45]), .CO(n94), .S(n95) );
  ADDFXL U148 ( .A(b[47]), .B(b[50]), .CI(b[48]), .CO(n88), .S(n89) );
  ADDFXL U149 ( .A(b[50]), .B(b[53]), .CI(b[51]), .CO(n82), .S(n83) );
  ADDFXL U150 ( .A(b[24]), .B(b[27]), .CI(b[25]), .CO(n134), .S(n135) );
  ADDFXL U151 ( .A(b[59]), .B(b[62]), .CI(b[60]), .CO(n64), .S(n65) );
  ADDFXL U152 ( .A(b[28]), .B(b[31]), .CI(b[29]), .CO(n126), .S(n127) );
  ADDFXL U153 ( .A(b[40]), .B(b[43]), .CI(b[41]), .CO(n102), .S(n103) );
  ADDFXL U154 ( .A(b[56]), .B(b[59]), .CI(b[57]), .CO(n70), .S(n71) );
  ADDFXL U155 ( .A(b[53]), .B(b[56]), .CI(b[54]), .CO(n76), .S(n77) );
  ADDHXL U156 ( .A(\b[0] ), .B(b[2]), .CO(n62), .S(product[2]) );
  ADDFXL U157 ( .A(n179), .B(n180), .CI(n60), .CO(n59), .S(product[5]) );
  ADDFXL U158 ( .A(n175), .B(n176), .CI(n58), .CO(n57), .S(product[7]) );
  ADDFXL U159 ( .A(n171), .B(n172), .CI(n56), .CO(n55), .S(product[9]) );
  ADDFXL U160 ( .A(n167), .B(n168), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U161 ( .A(n163), .B(n164), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U162 ( .A(n159), .B(n160), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U163 ( .A(n157), .B(n158), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U164 ( .A(n155), .B(n156), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U165 ( .A(n153), .B(n154), .CI(n47), .CO(n46), .S(product[18]) );
  ADDFXL U166 ( .A(n151), .B(n152), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U167 ( .A(n147), .B(n148), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U168 ( .A(n145), .B(n146), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U169 ( .A(n143), .B(n144), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U170 ( .A(n141), .B(n142), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U171 ( .A(n139), .B(n140), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U172 ( .A(n137), .B(n138), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U173 ( .A(n135), .B(n136), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U174 ( .A(n131), .B(n132), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U175 ( .A(n129), .B(n130), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U176 ( .A(n127), .B(n128), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U177 ( .A(n125), .B(n126), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U178 ( .A(n123), .B(n124), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U179 ( .A(n119), .B(n120), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U180 ( .A(n115), .B(n116), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U181 ( .A(n111), .B(n112), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U182 ( .A(n107), .B(n108), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U183 ( .A(n103), .B(n104), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U184 ( .A(n99), .B(n100), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U185 ( .A(n95), .B(n96), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U186 ( .A(n91), .B(n92), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U187 ( .A(n87), .B(n88), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U188 ( .A(n83), .B(n84), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U189 ( .A(n73), .B(n74), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U190 ( .A(n79), .B(n80), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U191 ( .A(n77), .B(n78), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U192 ( .A(n75), .B(n76), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U193 ( .A(n65), .B(n66), .CI(n3), .CO(n2), .S(product[62]) );
  ADDFXL U194 ( .A(n69), .B(n70), .CI(n5), .CO(n4), .S(product[60]) );
  XOR2X1 U195 ( .A(n323), .B(b[63]), .Y(n321) );
  ADDFXL U196 ( .A(n149), .B(n150), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U197 ( .A(n133), .B(n134), .CI(n37), .CO(n36), .S(product[28]) );
  ADDFXL U198 ( .A(n71), .B(n72), .CI(n6), .CO(n5), .S(product[59]) );
  XNOR2XL U199 ( .A(b[61]), .B(b[60]), .Y(n322) );
  ADDFXL U200 ( .A(n177), .B(n178), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U201 ( .A(n117), .B(n118), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U202 ( .A(n97), .B(n98), .CI(n19), .CO(n18), .S(product[46]) );
  XOR2X1 U203 ( .A(n321), .B(n322), .Y(product[63]) );
  XNOR2X1 U204 ( .A(n64), .B(n2), .Y(n323) );
endmodule


module GSIM_DW_mult_tc_4 ( a, b, product );
  input [3:0] a;
  input [63:0] b;
  output [67:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, \b[0] , \b[1] , n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318;
  assign product[1] = \b[0] ;
  assign \b[0]  = b[0];
  assign product[2] = \b[1] ;
  assign \b[1]  = b[1];

  ADDFXL U4 ( .A(b[60]), .B(n316), .CI(n4), .CO(n3), .S(product[61]) );
  ADDFXL U5 ( .A(b[59]), .B(n315), .CI(n5), .CO(n4), .S(product[60]) );
  ADDFXL U6 ( .A(b[58]), .B(n314), .CI(n6), .CO(n5), .S(product[59]) );
  ADDFXL U7 ( .A(b[57]), .B(n313), .CI(n7), .CO(n6), .S(product[58]) );
  ADDFXL U8 ( .A(b[56]), .B(n312), .CI(n8), .CO(n7), .S(product[57]) );
  ADDFXL U9 ( .A(b[55]), .B(n311), .CI(n9), .CO(n8), .S(product[56]) );
  ADDFXL U10 ( .A(b[54]), .B(n310), .CI(n10), .CO(n9), .S(product[55]) );
  ADDFXL U11 ( .A(b[53]), .B(n309), .CI(n11), .CO(n10), .S(product[54]) );
  ADDFXL U12 ( .A(b[52]), .B(n308), .CI(n12), .CO(n11), .S(product[53]) );
  ADDFXL U13 ( .A(b[51]), .B(n307), .CI(n13), .CO(n12), .S(product[52]) );
  ADDFXL U14 ( .A(b[50]), .B(n306), .CI(n14), .CO(n13), .S(product[51]) );
  ADDFXL U15 ( .A(b[49]), .B(n305), .CI(n15), .CO(n14), .S(product[50]) );
  ADDFXL U19 ( .A(b[45]), .B(n301), .CI(n19), .CO(n18), .S(product[46]) );
  ADDFXL U20 ( .A(b[44]), .B(n300), .CI(n20), .CO(n19), .S(product[45]) );
  ADDFXL U21 ( .A(b[43]), .B(n299), .CI(n21), .CO(n20), .S(product[44]) );
  ADDFXL U22 ( .A(b[42]), .B(n298), .CI(n22), .CO(n21), .S(product[43]) );
  ADDFXL U23 ( .A(b[41]), .B(n297), .CI(n23), .CO(n22), .S(product[42]) );
  ADDFXL U24 ( .A(b[40]), .B(n296), .CI(n24), .CO(n23), .S(product[41]) );
  ADDFXL U25 ( .A(b[39]), .B(n295), .CI(n25), .CO(n24), .S(product[40]) );
  ADDFXL U29 ( .A(b[35]), .B(n291), .CI(n29), .CO(n28), .S(product[36]) );
  ADDFXL U30 ( .A(b[34]), .B(n290), .CI(n30), .CO(n29), .S(product[35]) );
  ADDFXL U31 ( .A(b[33]), .B(n289), .CI(n31), .CO(n30), .S(product[34]) );
  ADDFXL U32 ( .A(b[32]), .B(n288), .CI(n32), .CO(n31), .S(product[33]) );
  ADDFXL U33 ( .A(b[31]), .B(n287), .CI(n33), .CO(n32), .S(product[32]) );
  ADDFXL U34 ( .A(b[30]), .B(n286), .CI(n34), .CO(n33), .S(product[31]) );
  ADDFXL U35 ( .A(b[29]), .B(n285), .CI(n35), .CO(n34), .S(product[30]) );
  ADDFXL U39 ( .A(b[25]), .B(n281), .CI(n39), .CO(n38), .S(product[26]) );
  ADDFXL U40 ( .A(b[24]), .B(n280), .CI(n40), .CO(n39), .S(product[25]) );
  ADDFXL U41 ( .A(b[23]), .B(n279), .CI(n41), .CO(n40), .S(product[24]) );
  ADDFXL U42 ( .A(b[22]), .B(n278), .CI(n42), .CO(n41), .S(product[23]) );
  ADDFXL U43 ( .A(b[21]), .B(n277), .CI(n43), .CO(n42), .S(product[22]) );
  ADDFXL U44 ( .A(b[20]), .B(n276), .CI(n44), .CO(n43), .S(product[21]) );
  ADDFXL U45 ( .A(b[19]), .B(n275), .CI(n45), .CO(n44), .S(product[20]) );
  ADDFXL U49 ( .A(b[15]), .B(n271), .CI(n49), .CO(n48), .S(product[16]) );
  ADDFXL U50 ( .A(b[14]), .B(n270), .CI(n50), .CO(n49), .S(product[15]) );
  ADDFXL U51 ( .A(b[13]), .B(n269), .CI(n51), .CO(n50), .S(product[14]) );
  ADDFXL U52 ( .A(b[12]), .B(n268), .CI(n52), .CO(n51), .S(product[13]) );
  ADDFXL U53 ( .A(b[11]), .B(n267), .CI(n53), .CO(n52), .S(product[12]) );
  ADDFXL U54 ( .A(b[10]), .B(n266), .CI(n54), .CO(n53), .S(product[11]) );
  ADDFXL U55 ( .A(b[9]), .B(n265), .CI(n55), .CO(n54), .S(product[10]) );
  ADDFXL U59 ( .A(b[5]), .B(n261), .CI(n59), .CO(n58), .S(product[6]) );
  ADDFXL U60 ( .A(b[4]), .B(n260), .CI(n60), .CO(n59), .S(product[5]) );
  CLKINVX6 U131 ( .A(b[2]), .Y(n260) );
  INVX1 U132 ( .A(\b[1] ), .Y(n259) );
  CLKINVX1 U133 ( .A(b[3]), .Y(n261) );
  ADDFHX1 U134 ( .A(b[3]), .B(n259), .CI(n61), .CO(n60), .S(product[4]) );
  XOR2XL U135 ( .A(b[2]), .B(\b[0] ), .Y(product[3]) );
  ADDFXL U136 ( .A(b[16]), .B(n272), .CI(n48), .CO(n47), .S(product[17]) );
  ADDFXL U137 ( .A(b[18]), .B(n274), .CI(n46), .CO(n45), .S(product[19]) );
  ADDFXL U138 ( .A(b[26]), .B(n282), .CI(n38), .CO(n37), .S(product[27]) );
  ADDFXL U139 ( .A(b[48]), .B(n304), .CI(n16), .CO(n15), .S(product[49]) );
  ADDFXL U140 ( .A(b[28]), .B(n284), .CI(n36), .CO(n35), .S(product[29]) );
  ADDFXL U141 ( .A(b[36]), .B(n292), .CI(n28), .CO(n27), .S(product[37]) );
  ADDFXL U142 ( .A(b[38]), .B(n294), .CI(n26), .CO(n25), .S(product[39]) );
  ADDFXL U143 ( .A(b[46]), .B(n302), .CI(n18), .CO(n17), .S(product[47]) );
  ADDFXL U144 ( .A(b[61]), .B(n317), .CI(n3), .CO(n2), .S(product[62]) );
  NAND2XL U145 ( .A(\b[0] ), .B(n260), .Y(n61) );
  INVXL U146 ( .A(b[20]), .Y(n278) );
  INVXL U147 ( .A(b[12]), .Y(n270) );
  INVXL U148 ( .A(b[13]), .Y(n271) );
  INVXL U149 ( .A(b[18]), .Y(n276) );
  INVXL U150 ( .A(b[10]), .Y(n268) );
  INVXL U151 ( .A(b[17]), .Y(n275) );
  INVXL U152 ( .A(b[19]), .Y(n277) );
  INVXL U153 ( .A(b[7]), .Y(n265) );
  INVXL U154 ( .A(b[8]), .Y(n266) );
  INVXL U155 ( .A(b[9]), .Y(n267) );
  INVXL U156 ( .A(b[11]), .Y(n269) );
  ADDFXL U157 ( .A(b[6]), .B(n262), .CI(n58), .CO(n57), .S(product[7]) );
  INVXL U158 ( .A(b[4]), .Y(n262) );
  INVXL U159 ( .A(b[14]), .Y(n272) );
  ADDFXL U160 ( .A(b[7]), .B(n263), .CI(n57), .CO(n56), .S(product[8]) );
  INVXL U161 ( .A(b[5]), .Y(n263) );
  ADDFXL U162 ( .A(b[8]), .B(n264), .CI(n56), .CO(n55), .S(product[9]) );
  INVXL U163 ( .A(b[6]), .Y(n264) );
  ADDFXL U164 ( .A(b[17]), .B(n273), .CI(n47), .CO(n46), .S(product[18]) );
  INVXL U165 ( .A(b[15]), .Y(n273) );
  INVXL U166 ( .A(b[16]), .Y(n274) );
  INVXL U167 ( .A(b[23]), .Y(n281) );
  INVXL U168 ( .A(b[58]), .Y(n316) );
  INVXL U169 ( .A(b[33]), .Y(n291) );
  INVXL U170 ( .A(b[43]), .Y(n301) );
  INVXL U171 ( .A(b[28]), .Y(n286) );
  INVXL U172 ( .A(b[38]), .Y(n296) );
  INVXL U173 ( .A(b[48]), .Y(n306) );
  INVXL U174 ( .A(b[27]), .Y(n285) );
  INVXL U175 ( .A(b[29]), .Y(n287) );
  INVXL U176 ( .A(b[30]), .Y(n288) );
  INVXL U177 ( .A(b[37]), .Y(n295) );
  INVXL U178 ( .A(b[39]), .Y(n297) );
  INVXL U179 ( .A(b[40]), .Y(n298) );
  INVXL U180 ( .A(b[47]), .Y(n305) );
  INVXL U181 ( .A(b[49]), .Y(n307) );
  INVXL U182 ( .A(b[50]), .Y(n308) );
  INVXL U183 ( .A(b[51]), .Y(n309) );
  INVXL U184 ( .A(b[21]), .Y(n279) );
  INVXL U185 ( .A(b[22]), .Y(n280) );
  INVXL U186 ( .A(b[31]), .Y(n289) );
  INVXL U187 ( .A(b[32]), .Y(n290) );
  INVXL U188 ( .A(b[41]), .Y(n299) );
  INVXL U189 ( .A(b[42]), .Y(n300) );
  INVXL U190 ( .A(b[52]), .Y(n310) );
  INVXL U191 ( .A(b[53]), .Y(n311) );
  INVXL U192 ( .A(b[54]), .Y(n312) );
  INVXL U193 ( .A(b[55]), .Y(n313) );
  INVXL U194 ( .A(b[56]), .Y(n314) );
  INVXL U195 ( .A(b[57]), .Y(n315) );
  XOR2X1 U196 ( .A(n318), .B(b[60]), .Y(product[63]) );
  INVXL U197 ( .A(b[59]), .Y(n317) );
  INVXL U198 ( .A(b[24]), .Y(n282) );
  INVXL U199 ( .A(b[34]), .Y(n292) );
  INVXL U200 ( .A(b[44]), .Y(n302) );
  ADDFXL U201 ( .A(b[27]), .B(n283), .CI(n37), .CO(n36), .S(product[28]) );
  INVXL U202 ( .A(b[25]), .Y(n283) );
  ADDFXL U203 ( .A(b[37]), .B(n293), .CI(n27), .CO(n26), .S(product[38]) );
  INVXL U204 ( .A(b[35]), .Y(n293) );
  ADDFXL U205 ( .A(b[47]), .B(n303), .CI(n17), .CO(n16), .S(product[48]) );
  INVXL U206 ( .A(b[45]), .Y(n303) );
  INVXL U207 ( .A(b[26]), .Y(n284) );
  INVXL U208 ( .A(b[36]), .Y(n294) );
  INVXL U209 ( .A(b[46]), .Y(n304) );
  XNOR2X1 U210 ( .A(n2), .B(b[62]), .Y(n318) );
endmodule


module GSIM_DW01_add_479 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;
  assign SUM[15] = B[15];
  assign SUM[14] = B[14];
  assign SUM[13] = B[13];
  assign SUM[12] = B[12];
  assign SUM[11] = B[11];
  assign SUM[10] = B[10];
  assign SUM[9] = B[9];
  assign SUM[8] = B[8];
  assign SUM[7] = B[7];
  assign SUM[6] = B[6];
  assign SUM[5] = B[5];
  assign SUM[4] = B[4];
  assign SUM[3] = B[3];
  assign SUM[2] = B[2];
  assign SUM[1] = B[1];

  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(n1), .CO(carry[18]), .S(SUM[17]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  AND2X2 U1 ( .A(B[16]), .B(A[16]), .Y(n1) );
  XOR2XL U2 ( .A(B[16]), .B(A[16]), .Y(SUM[16]) );
endmodule


module GSIM_DW01_add_478 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;
  assign SUM[0] = B[0];

  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2XL U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module GSIM_DW01_add_477 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;

  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFXL U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  ADDFXL U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  ADDFXL U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  ADDFXL U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  ADDFXL U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  ADDFXL U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFXL U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  ADDFXL U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  ADDFXL U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  ADDFXL U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFXL U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  ADDFXL U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  ADDFXL U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  ADDFXL U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  ADDFXL U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  ADDFXL U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  ADDFXL U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  ADDFXL U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  ADDFXL U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  ADDFXL U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  ADDFXL U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  XOR3X1 U1_63 ( .A(A[63]), .B(B[63]), .C(carry[63]), .Y(SUM[63]) );
  ADDFHX1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XL U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module GSIM ( clk, reset, in_en, b_in, out_valid, x_out );
  input [15:0] b_in;
  output [31:0] x_out;
  input clk, reset, in_en;
  output out_valid;
  wire   N1757, N1758, N1759, N1760, N1761, N1762, N1763, N1764, N1773, N1774,
         N1775, N1776, N1777, N1778, N1779, N1780, N1781, N1782, N1783, N1784,
         N1785, N1786, N1787, N1788, N1789, N1790, N1791, N1792, N1793, N1794,
         N1795, N1796, N1797, N1798, N1799, N1800, N1801, N1802, N1803, N1804,
         N1805, N1806, N1807, N1808, N1809, N1810, N1811, N1812, N1813, N1814,
         N1815, N1816, N1817, N1818, N1819, N1820, N1821, N1822, N1823, N1824,
         N1825, N1826, N1827, N1828, N1829, N1830, N1831, N1832, N1833, N1834,
         N1835, N1836, N1837, \bArray[0][63] , \bArray[0][62] ,
         \bArray[0][61] , \bArray[0][60] , \bArray[0][59] , \bArray[0][58] ,
         \bArray[0][57] , \bArray[0][56] , \bArray[0][55] , \bArray[0][54] ,
         \bArray[0][53] , \bArray[0][52] , \bArray[0][51] , \bArray[0][50] ,
         \bArray[0][49] , \bArray[0][48] , \bArray[0][47] , \bArray[0][46] ,
         \bArray[0][45] , \bArray[0][44] , \bArray[0][43] , \bArray[0][42] ,
         \bArray[0][41] , \bArray[0][40] , \bArray[0][39] , \bArray[0][38] ,
         \bArray[0][37] , \bArray[0][36] , \bArray[0][35] , \bArray[0][34] ,
         \bArray[0][33] , \bArray[0][32] , \bArray[0][31] , \bArray[0][30] ,
         \bArray[0][29] , \bArray[0][28] , \bArray[0][27] , \bArray[0][26] ,
         \bArray[0][25] , \bArray[0][24] , \bArray[0][23] , \bArray[0][22] ,
         \bArray[0][21] , \bArray[0][20] , \bArray[0][19] , \bArray[0][18] ,
         \bArray[0][17] , \bArray[0][16] , \bArray[1][63] , \bArray[1][62] ,
         \bArray[1][61] , \bArray[1][60] , \bArray[1][59] , \bArray[1][58] ,
         \bArray[1][57] , \bArray[1][56] , \bArray[1][55] , \bArray[1][54] ,
         \bArray[1][53] , \bArray[1][52] , \bArray[1][51] , \bArray[1][50] ,
         \bArray[1][49] , \bArray[1][48] , \bArray[1][47] , \bArray[1][46] ,
         \bArray[1][45] , \bArray[1][44] , \bArray[1][43] , \bArray[1][42] ,
         \bArray[1][41] , \bArray[1][40] , \bArray[1][39] , \bArray[1][38] ,
         \bArray[1][37] , \bArray[1][36] , \bArray[1][35] , \bArray[1][34] ,
         \bArray[1][33] , \bArray[1][32] , \bArray[1][31] , \bArray[1][30] ,
         \bArray[1][29] , \bArray[1][28] , \bArray[1][27] , \bArray[1][26] ,
         \bArray[1][25] , \bArray[1][24] , \bArray[1][23] , \bArray[1][22] ,
         \bArray[1][21] , \bArray[1][20] , \bArray[1][19] , \bArray[1][18] ,
         \bArray[1][17] , \bArray[1][16] , \bArray[2][63] , \bArray[2][62] ,
         \bArray[2][61] , \bArray[2][60] , \bArray[2][59] , \bArray[2][58] ,
         \bArray[2][57] , \bArray[2][56] , \bArray[2][55] , \bArray[2][54] ,
         \bArray[2][53] , \bArray[2][52] , \bArray[2][51] , \bArray[2][50] ,
         \bArray[2][49] , \bArray[2][48] , \bArray[2][47] , \bArray[2][46] ,
         \bArray[2][45] , \bArray[2][44] , \bArray[2][43] , \bArray[2][42] ,
         \bArray[2][41] , \bArray[2][40] , \bArray[2][39] , \bArray[2][38] ,
         \bArray[2][37] , \bArray[2][36] , \bArray[2][35] , \bArray[2][34] ,
         \bArray[2][33] , \bArray[2][32] , \bArray[2][31] , \bArray[2][30] ,
         \bArray[2][29] , \bArray[2][28] , \bArray[2][27] , \bArray[2][26] ,
         \bArray[2][25] , \bArray[2][24] , \bArray[2][23] , \bArray[2][22] ,
         \bArray[2][21] , \bArray[2][20] , \bArray[2][19] , \bArray[2][18] ,
         \bArray[2][17] , \bArray[2][16] , \bArray[3][63] , \bArray[3][62] ,
         \bArray[3][61] , \bArray[3][60] , \bArray[3][59] , \bArray[3][58] ,
         \bArray[3][57] , \bArray[3][56] , \bArray[3][55] , \bArray[3][54] ,
         \bArray[3][53] , \bArray[3][52] , \bArray[3][51] , \bArray[3][50] ,
         \bArray[3][49] , \bArray[3][48] , \bArray[3][47] , \bArray[3][46] ,
         \bArray[3][45] , \bArray[3][44] , \bArray[3][43] , \bArray[3][42] ,
         \bArray[3][41] , \bArray[3][40] , \bArray[3][39] , \bArray[3][38] ,
         \bArray[3][37] , \bArray[3][36] , \bArray[3][35] , \bArray[3][34] ,
         \bArray[3][33] , \bArray[3][32] , \bArray[3][31] , \bArray[3][30] ,
         \bArray[3][29] , \bArray[3][28] , \bArray[3][27] , \bArray[3][26] ,
         \bArray[3][25] , \bArray[3][24] , \bArray[3][23] , \bArray[3][22] ,
         \bArray[3][21] , \bArray[3][20] , \bArray[3][19] , \bArray[3][18] ,
         \bArray[3][17] , \bArray[3][16] , \bArray[4][63] , \bArray[4][62] ,
         \bArray[4][61] , \bArray[4][60] , \bArray[4][59] , \bArray[4][58] ,
         \bArray[4][57] , \bArray[4][56] , \bArray[4][55] , \bArray[4][54] ,
         \bArray[4][53] , \bArray[4][52] , \bArray[4][51] , \bArray[4][50] ,
         \bArray[4][49] , \bArray[4][48] , \bArray[4][47] , \bArray[4][46] ,
         \bArray[4][45] , \bArray[4][44] , \bArray[4][43] , \bArray[4][42] ,
         \bArray[4][41] , \bArray[4][40] , \bArray[4][39] , \bArray[4][38] ,
         \bArray[4][37] , \bArray[4][36] , \bArray[4][35] , \bArray[4][34] ,
         \bArray[4][33] , \bArray[4][32] , \bArray[4][31] , \bArray[4][30] ,
         \bArray[4][29] , \bArray[4][28] , \bArray[4][27] , \bArray[4][26] ,
         \bArray[4][25] , \bArray[4][24] , \bArray[4][23] , \bArray[4][22] ,
         \bArray[4][21] , \bArray[4][20] , \bArray[4][19] , \bArray[4][18] ,
         \bArray[4][17] , \bArray[4][16] , \bArray[5][63] , \bArray[5][62] ,
         \bArray[5][61] , \bArray[5][60] , \bArray[5][59] , \bArray[5][58] ,
         \bArray[5][57] , \bArray[5][56] , \bArray[5][55] , \bArray[5][54] ,
         \bArray[5][53] , \bArray[5][52] , \bArray[5][51] , \bArray[5][50] ,
         \bArray[5][49] , \bArray[5][48] , \bArray[5][47] , \bArray[5][46] ,
         \bArray[5][45] , \bArray[5][44] , \bArray[5][43] , \bArray[5][42] ,
         \bArray[5][41] , \bArray[5][40] , \bArray[5][39] , \bArray[5][38] ,
         \bArray[5][37] , \bArray[5][36] , \bArray[5][35] , \bArray[5][34] ,
         \bArray[5][33] , \bArray[5][32] , \bArray[5][31] , \bArray[5][30] ,
         \bArray[5][29] , \bArray[5][28] , \bArray[5][27] , \bArray[5][26] ,
         \bArray[5][25] , \bArray[5][24] , \bArray[5][23] , \bArray[5][22] ,
         \bArray[5][21] , \bArray[5][20] , \bArray[5][19] , \bArray[5][18] ,
         \bArray[5][17] , \bArray[5][16] , \bArray[6][63] , \bArray[6][62] ,
         \bArray[6][61] , \bArray[6][60] , \bArray[6][59] , \bArray[6][58] ,
         \bArray[6][57] , \bArray[6][56] , \bArray[6][55] , \bArray[6][54] ,
         \bArray[6][53] , \bArray[6][52] , \bArray[6][51] , \bArray[6][50] ,
         \bArray[6][49] , \bArray[6][48] , \bArray[6][47] , \bArray[6][46] ,
         \bArray[6][45] , \bArray[6][44] , \bArray[6][43] , \bArray[6][42] ,
         \bArray[6][41] , \bArray[6][40] , \bArray[6][39] , \bArray[6][38] ,
         \bArray[6][37] , \bArray[6][36] , \bArray[6][35] , \bArray[6][34] ,
         \bArray[6][33] , \bArray[6][32] , \bArray[6][31] , \bArray[6][30] ,
         \bArray[6][29] , \bArray[6][28] , \bArray[6][27] , \bArray[6][26] ,
         \bArray[6][25] , \bArray[6][24] , \bArray[6][23] , \bArray[6][22] ,
         \bArray[6][21] , \bArray[6][20] , \bArray[6][19] , \bArray[6][18] ,
         \bArray[6][17] , \bArray[6][16] , \bArray[7][63] , \bArray[7][62] ,
         \bArray[7][61] , \bArray[7][60] , \bArray[7][59] , \bArray[7][58] ,
         \bArray[7][57] , \bArray[7][56] , \bArray[7][55] , \bArray[7][54] ,
         \bArray[7][53] , \bArray[7][52] , \bArray[7][51] , \bArray[7][50] ,
         \bArray[7][49] , \bArray[7][48] , \bArray[7][47] , \bArray[7][46] ,
         \bArray[7][45] , \bArray[7][44] , \bArray[7][43] , \bArray[7][42] ,
         \bArray[7][41] , \bArray[7][40] , \bArray[7][39] , \bArray[7][38] ,
         \bArray[7][37] , \bArray[7][36] , \bArray[7][35] , \bArray[7][34] ,
         \bArray[7][33] , \bArray[7][32] , \bArray[7][31] , \bArray[7][30] ,
         \bArray[7][29] , \bArray[7][28] , \bArray[7][27] , \bArray[7][26] ,
         \bArray[7][25] , \bArray[7][24] , \bArray[7][23] , \bArray[7][22] ,
         \bArray[7][21] , \bArray[7][20] , \bArray[7][19] , \bArray[7][18] ,
         \bArray[7][17] , \bArray[7][16] , \bArray[8][63] , \bArray[8][62] ,
         \bArray[8][61] , \bArray[8][60] , \bArray[8][59] , \bArray[8][58] ,
         \bArray[8][57] , \bArray[8][56] , \bArray[8][55] , \bArray[8][54] ,
         \bArray[8][53] , \bArray[8][52] , \bArray[8][51] , \bArray[8][50] ,
         \bArray[8][49] , \bArray[8][48] , \bArray[8][47] , \bArray[8][46] ,
         \bArray[8][45] , \bArray[8][44] , \bArray[8][43] , \bArray[8][42] ,
         \bArray[8][41] , \bArray[8][40] , \bArray[8][39] , \bArray[8][38] ,
         \bArray[8][37] , \bArray[8][36] , \bArray[8][35] , \bArray[8][34] ,
         \bArray[8][33] , \bArray[8][32] , \bArray[8][31] , \bArray[8][30] ,
         \bArray[8][29] , \bArray[8][28] , \bArray[8][27] , \bArray[8][26] ,
         \bArray[8][25] , \bArray[8][24] , \bArray[8][23] , \bArray[8][22] ,
         \bArray[8][21] , \bArray[8][20] , \bArray[8][19] , \bArray[8][18] ,
         \bArray[8][17] , \bArray[8][16] , \bArray[9][63] , \bArray[9][62] ,
         \bArray[9][61] , \bArray[9][60] , \bArray[9][59] , \bArray[9][58] ,
         \bArray[9][57] , \bArray[9][56] , \bArray[9][55] , \bArray[9][54] ,
         \bArray[9][53] , \bArray[9][52] , \bArray[9][51] , \bArray[9][50] ,
         \bArray[9][49] , \bArray[9][48] , \bArray[9][47] , \bArray[9][46] ,
         \bArray[9][45] , \bArray[9][44] , \bArray[9][43] , \bArray[9][42] ,
         \bArray[9][41] , \bArray[9][40] , \bArray[9][39] , \bArray[9][38] ,
         \bArray[9][37] , \bArray[9][36] , \bArray[9][35] , \bArray[9][34] ,
         \bArray[9][33] , \bArray[9][32] , \bArray[9][31] , \bArray[9][30] ,
         \bArray[9][29] , \bArray[9][28] , \bArray[9][27] , \bArray[9][26] ,
         \bArray[9][25] , \bArray[9][24] , \bArray[9][23] , \bArray[9][22] ,
         \bArray[9][21] , \bArray[9][20] , \bArray[9][19] , \bArray[9][18] ,
         \bArray[9][17] , \bArray[9][16] , \bArray[10][63] , \bArray[10][62] ,
         \bArray[10][61] , \bArray[10][60] , \bArray[10][59] ,
         \bArray[10][58] , \bArray[10][57] , \bArray[10][56] ,
         \bArray[10][55] , \bArray[10][54] , \bArray[10][53] ,
         \bArray[10][52] , \bArray[10][51] , \bArray[10][50] ,
         \bArray[10][49] , \bArray[10][48] , \bArray[10][47] ,
         \bArray[10][46] , \bArray[10][45] , \bArray[10][44] ,
         \bArray[10][43] , \bArray[10][42] , \bArray[10][41] ,
         \bArray[10][40] , \bArray[10][39] , \bArray[10][38] ,
         \bArray[10][37] , \bArray[10][36] , \bArray[10][35] ,
         \bArray[10][34] , \bArray[10][33] , \bArray[10][32] ,
         \bArray[10][31] , \bArray[10][30] , \bArray[10][29] ,
         \bArray[10][28] , \bArray[10][27] , \bArray[10][26] ,
         \bArray[10][25] , \bArray[10][24] , \bArray[10][23] ,
         \bArray[10][22] , \bArray[10][21] , \bArray[10][20] ,
         \bArray[10][19] , \bArray[10][18] , \bArray[10][17] ,
         \bArray[10][16] , \bArray[11][63] , \bArray[11][62] ,
         \bArray[11][61] , \bArray[11][60] , \bArray[11][59] ,
         \bArray[11][58] , \bArray[11][57] , \bArray[11][56] ,
         \bArray[11][55] , \bArray[11][54] , \bArray[11][53] ,
         \bArray[11][52] , \bArray[11][51] , \bArray[11][50] ,
         \bArray[11][49] , \bArray[11][48] , \bArray[11][47] ,
         \bArray[11][46] , \bArray[11][45] , \bArray[11][44] ,
         \bArray[11][43] , \bArray[11][42] , \bArray[11][41] ,
         \bArray[11][40] , \bArray[11][39] , \bArray[11][38] ,
         \bArray[11][37] , \bArray[11][36] , \bArray[11][35] ,
         \bArray[11][34] , \bArray[11][33] , \bArray[11][32] ,
         \bArray[11][31] , \bArray[11][30] , \bArray[11][29] ,
         \bArray[11][28] , \bArray[11][27] , \bArray[11][26] ,
         \bArray[11][25] , \bArray[11][24] , \bArray[11][23] ,
         \bArray[11][22] , \bArray[11][21] , \bArray[11][20] ,
         \bArray[11][19] , \bArray[11][18] , \bArray[11][17] ,
         \bArray[11][16] , \bArray[12][63] , \bArray[12][62] ,
         \bArray[12][61] , \bArray[12][60] , \bArray[12][59] ,
         \bArray[12][58] , \bArray[12][57] , \bArray[12][56] ,
         \bArray[12][55] , \bArray[12][54] , \bArray[12][53] ,
         \bArray[12][52] , \bArray[12][51] , \bArray[12][50] ,
         \bArray[12][49] , \bArray[12][48] , \bArray[12][47] ,
         \bArray[12][46] , \bArray[12][45] , \bArray[12][44] ,
         \bArray[12][43] , \bArray[12][42] , \bArray[12][41] ,
         \bArray[12][40] , \bArray[12][39] , \bArray[12][38] ,
         \bArray[12][37] , \bArray[12][36] , \bArray[12][35] ,
         \bArray[12][34] , \bArray[12][33] , \bArray[12][32] ,
         \bArray[12][31] , \bArray[12][30] , \bArray[12][29] ,
         \bArray[12][28] , \bArray[12][27] , \bArray[12][26] ,
         \bArray[12][25] , \bArray[12][24] , \bArray[12][23] ,
         \bArray[12][22] , \bArray[12][21] , \bArray[12][20] ,
         \bArray[12][19] , \bArray[12][18] , \bArray[12][17] ,
         \bArray[12][16] , \bArray[13][63] , \bArray[13][62] ,
         \bArray[13][61] , \bArray[13][60] , \bArray[13][59] ,
         \bArray[13][58] , \bArray[13][57] , \bArray[13][56] ,
         \bArray[13][55] , \bArray[13][54] , \bArray[13][53] ,
         \bArray[13][52] , \bArray[13][51] , \bArray[13][50] ,
         \bArray[13][49] , \bArray[13][48] , \bArray[13][47] ,
         \bArray[13][46] , \bArray[13][45] , \bArray[13][44] ,
         \bArray[13][43] , \bArray[13][42] , \bArray[13][41] ,
         \bArray[13][40] , \bArray[13][39] , \bArray[13][38] ,
         \bArray[13][37] , \bArray[13][36] , \bArray[13][35] ,
         \bArray[13][34] , \bArray[13][33] , \bArray[13][32] ,
         \bArray[13][31] , \bArray[13][30] , \bArray[13][29] ,
         \bArray[13][28] , \bArray[13][27] , \bArray[13][26] ,
         \bArray[13][25] , \bArray[13][24] , \bArray[13][23] ,
         \bArray[13][22] , \bArray[13][21] , \bArray[13][20] ,
         \bArray[13][19] , \bArray[13][18] , \bArray[13][17] ,
         \bArray[13][16] , \bArray[14][63] , \bArray[14][62] ,
         \bArray[14][61] , \bArray[14][60] , \bArray[14][59] ,
         \bArray[14][58] , \bArray[14][57] , \bArray[14][56] ,
         \bArray[14][55] , \bArray[14][54] , \bArray[14][53] ,
         \bArray[14][52] , \bArray[14][51] , \bArray[14][50] ,
         \bArray[14][49] , \bArray[14][48] , \bArray[14][47] ,
         \bArray[14][46] , \bArray[14][45] , \bArray[14][44] ,
         \bArray[14][43] , \bArray[14][42] , \bArray[14][41] ,
         \bArray[14][40] , \bArray[14][39] , \bArray[14][38] ,
         \bArray[14][37] , \bArray[14][36] , \bArray[14][35] ,
         \bArray[14][34] , \bArray[14][33] , \bArray[14][32] ,
         \bArray[14][31] , \bArray[14][30] , \bArray[14][29] ,
         \bArray[14][28] , \bArray[14][27] , \bArray[14][26] ,
         \bArray[14][25] , \bArray[14][24] , \bArray[14][23] ,
         \bArray[14][22] , \bArray[14][21] , \bArray[14][20] ,
         \bArray[14][19] , \bArray[14][18] , \bArray[14][17] ,
         \bArray[14][16] , \bArray[15][63] , \bArray[15][62] ,
         \bArray[15][61] , \bArray[15][60] , \bArray[15][59] ,
         \bArray[15][58] , \bArray[15][57] , \bArray[15][56] ,
         \bArray[15][55] , \bArray[15][54] , \bArray[15][53] ,
         \bArray[15][52] , \bArray[15][51] , \bArray[15][50] ,
         \bArray[15][49] , \bArray[15][48] , \bArray[15][47] ,
         \bArray[15][46] , \bArray[15][45] , \bArray[15][44] ,
         \bArray[15][43] , \bArray[15][42] , \bArray[15][41] ,
         \bArray[15][40] , \bArray[15][39] , \bArray[15][38] ,
         \bArray[15][37] , \bArray[15][36] , \bArray[15][35] ,
         \bArray[15][34] , \bArray[15][33] , \bArray[15][32] ,
         \bArray[15][31] , \bArray[15][30] , \bArray[15][29] ,
         \bArray[15][28] , \bArray[15][27] , \bArray[15][26] ,
         \bArray[15][25] , \bArray[15][24] , \bArray[15][23] ,
         \bArray[15][22] , \bArray[15][21] , \bArray[15][20] ,
         \bArray[15][19] , \bArray[15][18] , \bArray[15][17] ,
         \bArray[15][16] , N2348, \xArray[0][63] , \xArray[0][62] ,
         \xArray[0][61] , \xArray[0][60] , \xArray[0][59] , \xArray[0][58] ,
         \xArray[0][57] , \xArray[0][56] , \xArray[0][55] , \xArray[0][54] ,
         \xArray[0][53] , \xArray[0][52] , \xArray[0][51] , \xArray[0][50] ,
         \xArray[0][49] , \xArray[0][48] , \xArray[0][47] , \xArray[0][46] ,
         \xArray[0][45] , \xArray[0][44] , \xArray[0][43] , \xArray[0][42] ,
         \xArray[0][41] , \xArray[0][40] , \xArray[0][39] , \xArray[0][38] ,
         \xArray[0][37] , \xArray[0][36] , \xArray[0][35] , \xArray[0][34] ,
         \xArray[0][33] , \xArray[0][32] , \xArray[0][31] , \xArray[0][30] ,
         \xArray[0][29] , \xArray[0][28] , \xArray[0][27] , \xArray[0][26] ,
         \xArray[0][25] , \xArray[0][24] , \xArray[0][23] , \xArray[0][22] ,
         \xArray[0][21] , \xArray[0][20] , \xArray[0][19] , \xArray[0][18] ,
         \xArray[0][17] , \xArray[0][16] , \xArray[0][15] , \xArray[0][14] ,
         \xArray[0][13] , \xArray[0][12] , \xArray[0][11] , \xArray[0][10] ,
         \xArray[0][9] , \xArray[0][8] , \xArray[0][7] , \xArray[0][6] ,
         \xArray[0][5] , \xArray[0][4] , \xArray[0][3] , \xArray[0][2] ,
         \xArray[0][1] , \xArray[0][0] , \xArray[1][63] , \xArray[1][62] ,
         \xArray[1][61] , \xArray[1][60] , \xArray[1][59] , \xArray[1][58] ,
         \xArray[1][57] , \xArray[1][56] , \xArray[1][55] , \xArray[1][54] ,
         \xArray[1][53] , \xArray[1][52] , \xArray[1][51] , \xArray[1][50] ,
         \xArray[1][49] , \xArray[1][48] , \xArray[1][47] , \xArray[1][46] ,
         \xArray[1][45] , \xArray[1][44] , \xArray[1][43] , \xArray[1][42] ,
         \xArray[1][41] , \xArray[1][40] , \xArray[1][39] , \xArray[1][38] ,
         \xArray[1][37] , \xArray[1][36] , \xArray[1][35] , \xArray[1][34] ,
         \xArray[1][33] , \xArray[1][32] , \xArray[1][31] , \xArray[1][30] ,
         \xArray[1][29] , \xArray[1][28] , \xArray[1][27] , \xArray[1][26] ,
         \xArray[1][25] , \xArray[1][24] , \xArray[1][23] , \xArray[1][22] ,
         \xArray[1][21] , \xArray[1][20] , \xArray[1][19] , \xArray[1][18] ,
         \xArray[1][17] , \xArray[1][16] , \xArray[1][15] , \xArray[1][14] ,
         \xArray[1][13] , \xArray[1][12] , \xArray[1][11] , \xArray[1][10] ,
         \xArray[1][9] , \xArray[1][8] , \xArray[1][7] , \xArray[1][6] ,
         \xArray[1][5] , \xArray[1][4] , \xArray[1][3] , \xArray[1][2] ,
         \xArray[1][1] , \xArray[1][0] , \xArray[2][63] , \xArray[2][62] ,
         \xArray[2][61] , \xArray[2][60] , \xArray[2][59] , \xArray[2][58] ,
         \xArray[2][57] , \xArray[2][56] , \xArray[2][55] , \xArray[2][54] ,
         \xArray[2][53] , \xArray[2][52] , \xArray[2][51] , \xArray[2][50] ,
         \xArray[2][49] , \xArray[2][48] , \xArray[2][47] , \xArray[2][46] ,
         \xArray[2][45] , \xArray[2][44] , \xArray[2][43] , \xArray[2][42] ,
         \xArray[2][41] , \xArray[2][40] , \xArray[2][39] , \xArray[2][38] ,
         \xArray[2][37] , \xArray[2][36] , \xArray[2][35] , \xArray[2][34] ,
         \xArray[2][33] , \xArray[2][32] , \xArray[2][31] , \xArray[2][30] ,
         \xArray[2][29] , \xArray[2][28] , \xArray[2][27] , \xArray[2][26] ,
         \xArray[2][25] , \xArray[2][24] , \xArray[2][23] , \xArray[2][22] ,
         \xArray[2][21] , \xArray[2][20] , \xArray[2][19] , \xArray[2][18] ,
         \xArray[2][17] , \xArray[2][16] , \xArray[2][15] , \xArray[2][14] ,
         \xArray[2][13] , \xArray[2][12] , \xArray[2][11] , \xArray[2][10] ,
         \xArray[2][9] , \xArray[2][8] , \xArray[2][7] , \xArray[2][6] ,
         \xArray[2][5] , \xArray[2][4] , \xArray[2][3] , \xArray[2][2] ,
         \xArray[2][1] , \xArray[2][0] , \xArray[3][63] , \xArray[3][62] ,
         \xArray[3][61] , \xArray[3][60] , \xArray[3][59] , \xArray[3][58] ,
         \xArray[3][57] , \xArray[3][56] , \xArray[3][55] , \xArray[3][54] ,
         \xArray[3][53] , \xArray[3][52] , \xArray[3][51] , \xArray[3][50] ,
         \xArray[3][49] , \xArray[3][48] , \xArray[3][47] , \xArray[3][46] ,
         \xArray[3][45] , \xArray[3][44] , \xArray[3][43] , \xArray[3][42] ,
         \xArray[3][41] , \xArray[3][40] , \xArray[3][39] , \xArray[3][38] ,
         \xArray[3][37] , \xArray[3][36] , \xArray[3][35] , \xArray[3][34] ,
         \xArray[3][33] , \xArray[3][32] , \xArray[3][31] , \xArray[3][30] ,
         \xArray[3][29] , \xArray[3][28] , \xArray[3][27] , \xArray[3][26] ,
         \xArray[3][25] , \xArray[3][24] , \xArray[3][23] , \xArray[3][22] ,
         \xArray[3][21] , \xArray[3][20] , \xArray[3][19] , \xArray[3][18] ,
         \xArray[3][17] , \xArray[3][16] , \xArray[3][15] , \xArray[3][14] ,
         \xArray[3][13] , \xArray[3][12] , \xArray[3][11] , \xArray[3][10] ,
         \xArray[3][9] , \xArray[3][8] , \xArray[3][7] , \xArray[3][6] ,
         \xArray[3][5] , \xArray[3][4] , \xArray[3][3] , \xArray[3][2] ,
         \xArray[3][1] , \xArray[3][0] , \xArray[4][63] , \xArray[4][62] ,
         \xArray[4][61] , \xArray[4][60] , \xArray[4][59] , \xArray[4][58] ,
         \xArray[4][57] , \xArray[4][56] , \xArray[4][55] , \xArray[4][54] ,
         \xArray[4][53] , \xArray[4][52] , \xArray[4][51] , \xArray[4][50] ,
         \xArray[4][49] , \xArray[4][48] , \xArray[4][47] , \xArray[4][46] ,
         \xArray[4][45] , \xArray[4][44] , \xArray[4][43] , \xArray[4][42] ,
         \xArray[4][41] , \xArray[4][40] , \xArray[4][39] , \xArray[4][38] ,
         \xArray[4][37] , \xArray[4][36] , \xArray[4][35] , \xArray[4][34] ,
         \xArray[4][33] , \xArray[4][32] , \xArray[4][31] , \xArray[4][30] ,
         \xArray[4][29] , \xArray[4][28] , \xArray[4][27] , \xArray[4][26] ,
         \xArray[4][25] , \xArray[4][24] , \xArray[4][23] , \xArray[4][22] ,
         \xArray[4][21] , \xArray[4][20] , \xArray[4][19] , \xArray[4][18] ,
         \xArray[4][17] , \xArray[4][16] , \xArray[4][15] , \xArray[4][14] ,
         \xArray[4][13] , \xArray[4][12] , \xArray[4][11] , \xArray[4][10] ,
         \xArray[4][9] , \xArray[4][8] , \xArray[4][7] , \xArray[4][6] ,
         \xArray[4][5] , \xArray[4][4] , \xArray[4][3] , \xArray[4][2] ,
         \xArray[4][1] , \xArray[4][0] , \xArray[5][63] , \xArray[5][62] ,
         \xArray[5][61] , \xArray[5][60] , \xArray[5][59] , \xArray[5][58] ,
         \xArray[5][57] , \xArray[5][56] , \xArray[5][55] , \xArray[5][54] ,
         \xArray[5][53] , \xArray[5][52] , \xArray[5][51] , \xArray[5][50] ,
         \xArray[5][49] , \xArray[5][48] , \xArray[5][47] , \xArray[5][46] ,
         \xArray[5][45] , \xArray[5][44] , \xArray[5][43] , \xArray[5][42] ,
         \xArray[5][41] , \xArray[5][40] , \xArray[5][39] , \xArray[5][38] ,
         \xArray[5][37] , \xArray[5][36] , \xArray[5][35] , \xArray[5][34] ,
         \xArray[5][33] , \xArray[5][32] , \xArray[5][31] , \xArray[5][30] ,
         \xArray[5][29] , \xArray[5][28] , \xArray[5][27] , \xArray[5][26] ,
         \xArray[5][25] , \xArray[5][24] , \xArray[5][23] , \xArray[5][22] ,
         \xArray[5][21] , \xArray[5][20] , \xArray[5][19] , \xArray[5][18] ,
         \xArray[5][17] , \xArray[5][16] , \xArray[5][15] , \xArray[5][14] ,
         \xArray[5][13] , \xArray[5][12] , \xArray[5][11] , \xArray[5][10] ,
         \xArray[5][9] , \xArray[5][8] , \xArray[5][7] , \xArray[5][6] ,
         \xArray[5][5] , \xArray[5][4] , \xArray[5][3] , \xArray[5][2] ,
         \xArray[5][1] , \xArray[5][0] , \xArray[6][63] , \xArray[6][62] ,
         \xArray[6][61] , \xArray[6][60] , \xArray[6][59] , \xArray[6][58] ,
         \xArray[6][57] , \xArray[6][56] , \xArray[6][55] , \xArray[6][54] ,
         \xArray[6][53] , \xArray[6][52] , \xArray[6][51] , \xArray[6][50] ,
         \xArray[6][49] , \xArray[6][48] , \xArray[6][47] , \xArray[6][46] ,
         \xArray[6][45] , \xArray[6][44] , \xArray[6][43] , \xArray[6][42] ,
         \xArray[6][41] , \xArray[6][40] , \xArray[6][39] , \xArray[6][38] ,
         \xArray[6][37] , \xArray[6][36] , \xArray[6][35] , \xArray[6][34] ,
         \xArray[6][33] , \xArray[6][32] , \xArray[6][31] , \xArray[6][30] ,
         \xArray[6][29] , \xArray[6][28] , \xArray[6][27] , \xArray[6][26] ,
         \xArray[6][25] , \xArray[6][24] , \xArray[6][23] , \xArray[6][22] ,
         \xArray[6][21] , \xArray[6][20] , \xArray[6][19] , \xArray[6][18] ,
         \xArray[6][17] , \xArray[6][16] , \xArray[6][15] , \xArray[6][14] ,
         \xArray[6][13] , \xArray[6][12] , \xArray[6][11] , \xArray[6][10] ,
         \xArray[6][9] , \xArray[6][8] , \xArray[6][7] , \xArray[6][6] ,
         \xArray[6][5] , \xArray[6][4] , \xArray[6][3] , \xArray[6][2] ,
         \xArray[6][1] , \xArray[6][0] , \xArray[7][63] , \xArray[7][62] ,
         \xArray[7][61] , \xArray[7][60] , \xArray[7][59] , \xArray[7][58] ,
         \xArray[7][57] , \xArray[7][56] , \xArray[7][55] , \xArray[7][54] ,
         \xArray[7][53] , \xArray[7][52] , \xArray[7][51] , \xArray[7][50] ,
         \xArray[7][49] , \xArray[7][48] , \xArray[7][47] , \xArray[7][46] ,
         \xArray[7][45] , \xArray[7][44] , \xArray[7][43] , \xArray[7][42] ,
         \xArray[7][41] , \xArray[7][40] , \xArray[7][39] , \xArray[7][38] ,
         \xArray[7][37] , \xArray[7][36] , \xArray[7][35] , \xArray[7][34] ,
         \xArray[7][33] , \xArray[7][32] , \xArray[7][31] , \xArray[7][30] ,
         \xArray[7][29] , \xArray[7][28] , \xArray[7][27] , \xArray[7][26] ,
         \xArray[7][25] , \xArray[7][24] , \xArray[7][23] , \xArray[7][22] ,
         \xArray[7][21] , \xArray[7][20] , \xArray[7][19] , \xArray[7][18] ,
         \xArray[7][17] , \xArray[7][16] , \xArray[7][15] , \xArray[7][14] ,
         \xArray[7][13] , \xArray[7][12] , \xArray[7][11] , \xArray[7][10] ,
         \xArray[7][9] , \xArray[7][8] , \xArray[7][7] , \xArray[7][6] ,
         \xArray[7][5] , \xArray[7][4] , \xArray[7][3] , \xArray[7][2] ,
         \xArray[7][1] , \xArray[7][0] , \xArray[8][63] , \xArray[8][62] ,
         \xArray[8][61] , \xArray[8][60] , \xArray[8][59] , \xArray[8][58] ,
         \xArray[8][57] , \xArray[8][56] , \xArray[8][55] , \xArray[8][54] ,
         \xArray[8][53] , \xArray[8][52] , \xArray[8][51] , \xArray[8][50] ,
         \xArray[8][49] , \xArray[8][48] , \xArray[8][47] , \xArray[8][46] ,
         \xArray[8][45] , \xArray[8][44] , \xArray[8][43] , \xArray[8][42] ,
         \xArray[8][41] , \xArray[8][40] , \xArray[8][39] , \xArray[8][38] ,
         \xArray[8][37] , \xArray[8][36] , \xArray[8][35] , \xArray[8][34] ,
         \xArray[8][33] , \xArray[8][32] , \xArray[8][31] , \xArray[8][30] ,
         \xArray[8][29] , \xArray[8][28] , \xArray[8][27] , \xArray[8][26] ,
         \xArray[8][25] , \xArray[8][24] , \xArray[8][23] , \xArray[8][22] ,
         \xArray[8][21] , \xArray[8][20] , \xArray[8][19] , \xArray[8][18] ,
         \xArray[8][17] , \xArray[8][16] , \xArray[8][15] , \xArray[8][14] ,
         \xArray[8][13] , \xArray[8][12] , \xArray[8][11] , \xArray[8][10] ,
         \xArray[8][9] , \xArray[8][8] , \xArray[8][7] , \xArray[8][6] ,
         \xArray[8][5] , \xArray[8][4] , \xArray[8][3] , \xArray[8][2] ,
         \xArray[8][1] , \xArray[8][0] , \xArray[9][63] , \xArray[9][62] ,
         \xArray[9][61] , \xArray[9][60] , \xArray[9][59] , \xArray[9][58] ,
         \xArray[9][57] , \xArray[9][56] , \xArray[9][55] , \xArray[9][54] ,
         \xArray[9][53] , \xArray[9][52] , \xArray[9][51] , \xArray[9][50] ,
         \xArray[9][49] , \xArray[9][48] , \xArray[9][47] , \xArray[9][46] ,
         \xArray[9][45] , \xArray[9][44] , \xArray[9][43] , \xArray[9][42] ,
         \xArray[9][41] , \xArray[9][40] , \xArray[9][39] , \xArray[9][38] ,
         \xArray[9][37] , \xArray[9][36] , \xArray[9][35] , \xArray[9][34] ,
         \xArray[9][33] , \xArray[9][32] , \xArray[9][31] , \xArray[9][30] ,
         \xArray[9][29] , \xArray[9][28] , \xArray[9][27] , \xArray[9][26] ,
         \xArray[9][25] , \xArray[9][24] , \xArray[9][23] , \xArray[9][22] ,
         \xArray[9][21] , \xArray[9][20] , \xArray[9][19] , \xArray[9][18] ,
         \xArray[9][17] , \xArray[9][16] , \xArray[9][15] , \xArray[9][14] ,
         \xArray[9][13] , \xArray[9][12] , \xArray[9][11] , \xArray[9][10] ,
         \xArray[9][9] , \xArray[9][8] , \xArray[9][7] , \xArray[9][6] ,
         \xArray[9][5] , \xArray[9][4] , \xArray[9][3] , \xArray[9][2] ,
         \xArray[9][1] , \xArray[9][0] , \xArray[10][63] , \xArray[10][62] ,
         \xArray[10][61] , \xArray[10][60] , \xArray[10][59] ,
         \xArray[10][58] , \xArray[10][57] , \xArray[10][56] ,
         \xArray[10][55] , \xArray[10][54] , \xArray[10][53] ,
         \xArray[10][52] , \xArray[10][51] , \xArray[10][50] ,
         \xArray[10][49] , \xArray[10][48] , \xArray[10][47] ,
         \xArray[10][46] , \xArray[10][45] , \xArray[10][44] ,
         \xArray[10][43] , \xArray[10][42] , \xArray[10][41] ,
         \xArray[10][40] , \xArray[10][39] , \xArray[10][38] ,
         \xArray[10][37] , \xArray[10][36] , \xArray[10][35] ,
         \xArray[10][34] , \xArray[10][33] , \xArray[10][32] ,
         \xArray[10][31] , \xArray[10][30] , \xArray[10][29] ,
         \xArray[10][28] , \xArray[10][27] , \xArray[10][26] ,
         \xArray[10][25] , \xArray[10][24] , \xArray[10][23] ,
         \xArray[10][22] , \xArray[10][21] , \xArray[10][20] ,
         \xArray[10][19] , \xArray[10][18] , \xArray[10][17] ,
         \xArray[10][16] , \xArray[10][15] , \xArray[10][14] ,
         \xArray[10][13] , \xArray[10][12] , \xArray[10][11] ,
         \xArray[10][10] , \xArray[10][9] , \xArray[10][8] , \xArray[10][7] ,
         \xArray[10][6] , \xArray[10][5] , \xArray[10][4] , \xArray[10][3] ,
         \xArray[10][2] , \xArray[10][1] , \xArray[10][0] , \xArray[11][63] ,
         \xArray[11][62] , \xArray[11][61] , \xArray[11][60] ,
         \xArray[11][59] , \xArray[11][58] , \xArray[11][57] ,
         \xArray[11][56] , \xArray[11][55] , \xArray[11][54] ,
         \xArray[11][53] , \xArray[11][52] , \xArray[11][51] ,
         \xArray[11][50] , \xArray[11][49] , \xArray[11][48] ,
         \xArray[11][47] , \xArray[11][46] , \xArray[11][45] ,
         \xArray[11][44] , \xArray[11][43] , \xArray[11][42] ,
         \xArray[11][41] , \xArray[11][40] , \xArray[11][39] ,
         \xArray[11][38] , \xArray[11][37] , \xArray[11][36] ,
         \xArray[11][35] , \xArray[11][34] , \xArray[11][33] ,
         \xArray[11][32] , \xArray[11][31] , \xArray[11][30] ,
         \xArray[11][29] , \xArray[11][28] , \xArray[11][27] ,
         \xArray[11][26] , \xArray[11][25] , \xArray[11][24] ,
         \xArray[11][23] , \xArray[11][22] , \xArray[11][21] ,
         \xArray[11][20] , \xArray[11][19] , \xArray[11][18] ,
         \xArray[11][17] , \xArray[11][16] , \xArray[11][15] ,
         \xArray[11][14] , \xArray[11][13] , \xArray[11][12] ,
         \xArray[11][11] , \xArray[11][10] , \xArray[11][9] , \xArray[11][8] ,
         \xArray[11][7] , \xArray[11][6] , \xArray[11][5] , \xArray[11][4] ,
         \xArray[11][3] , \xArray[11][2] , \xArray[11][1] , \xArray[11][0] ,
         \xArray[12][63] , \xArray[12][62] , \xArray[12][61] ,
         \xArray[12][60] , \xArray[12][59] , \xArray[12][58] ,
         \xArray[12][57] , \xArray[12][56] , \xArray[12][55] ,
         \xArray[12][54] , \xArray[12][53] , \xArray[12][52] ,
         \xArray[12][51] , \xArray[12][50] , \xArray[12][49] ,
         \xArray[12][48] , \xArray[12][47] , \xArray[12][46] ,
         \xArray[12][45] , \xArray[12][44] , \xArray[12][43] ,
         \xArray[12][42] , \xArray[12][41] , \xArray[12][40] ,
         \xArray[12][39] , \xArray[12][38] , \xArray[12][37] ,
         \xArray[12][36] , \xArray[12][35] , \xArray[12][34] ,
         \xArray[12][33] , \xArray[12][32] , \xArray[12][31] ,
         \xArray[12][30] , \xArray[12][29] , \xArray[12][28] ,
         \xArray[12][27] , \xArray[12][26] , \xArray[12][25] ,
         \xArray[12][24] , \xArray[12][23] , \xArray[12][22] ,
         \xArray[12][21] , \xArray[12][20] , \xArray[12][19] ,
         \xArray[12][18] , \xArray[12][17] , \xArray[12][16] ,
         \xArray[12][15] , \xArray[12][14] , \xArray[12][13] ,
         \xArray[12][12] , \xArray[12][11] , \xArray[12][10] , \xArray[12][9] ,
         \xArray[12][8] , \xArray[12][7] , \xArray[12][6] , \xArray[12][5] ,
         \xArray[12][4] , \xArray[12][3] , \xArray[12][2] , \xArray[12][1] ,
         \xArray[12][0] , \xArray[13][63] , \xArray[13][62] , \xArray[13][61] ,
         \xArray[13][60] , \xArray[13][59] , \xArray[13][58] ,
         \xArray[13][57] , \xArray[13][56] , \xArray[13][55] ,
         \xArray[13][54] , \xArray[13][53] , \xArray[13][52] ,
         \xArray[13][51] , \xArray[13][50] , \xArray[13][49] ,
         \xArray[13][48] , \xArray[13][47] , \xArray[13][46] ,
         \xArray[13][45] , \xArray[13][44] , \xArray[13][43] ,
         \xArray[13][42] , \xArray[13][41] , \xArray[13][40] ,
         \xArray[13][39] , \xArray[13][38] , \xArray[13][37] ,
         \xArray[13][36] , \xArray[13][35] , \xArray[13][34] ,
         \xArray[13][33] , \xArray[13][32] , \xArray[13][31] ,
         \xArray[13][30] , \xArray[13][29] , \xArray[13][28] ,
         \xArray[13][27] , \xArray[13][26] , \xArray[13][25] ,
         \xArray[13][24] , \xArray[13][23] , \xArray[13][22] ,
         \xArray[13][21] , \xArray[13][20] , \xArray[13][19] ,
         \xArray[13][18] , \xArray[13][17] , \xArray[13][16] ,
         \xArray[13][15] , \xArray[13][14] , \xArray[13][13] ,
         \xArray[13][12] , \xArray[13][11] , \xArray[13][10] , \xArray[13][9] ,
         \xArray[13][8] , \xArray[13][7] , \xArray[13][6] , \xArray[13][5] ,
         \xArray[13][4] , \xArray[13][3] , \xArray[13][2] , \xArray[13][1] ,
         \xArray[13][0] , \xArray[14][63] , \xArray[14][62] , \xArray[14][61] ,
         \xArray[14][60] , \xArray[14][59] , \xArray[14][58] ,
         \xArray[14][57] , \xArray[14][56] , \xArray[14][55] ,
         \xArray[14][54] , \xArray[14][53] , \xArray[14][52] ,
         \xArray[14][51] , \xArray[14][50] , \xArray[14][49] ,
         \xArray[14][48] , \xArray[14][47] , \xArray[14][46] ,
         \xArray[14][45] , \xArray[14][44] , \xArray[14][43] ,
         \xArray[14][42] , \xArray[14][41] , \xArray[14][40] ,
         \xArray[14][39] , \xArray[14][38] , \xArray[14][37] ,
         \xArray[14][36] , \xArray[14][35] , \xArray[14][34] ,
         \xArray[14][33] , \xArray[14][32] , \xArray[14][31] ,
         \xArray[14][30] , \xArray[14][29] , \xArray[14][28] ,
         \xArray[14][27] , \xArray[14][26] , \xArray[14][25] ,
         \xArray[14][24] , \xArray[14][23] , \xArray[14][22] ,
         \xArray[14][21] , \xArray[14][20] , \xArray[14][19] ,
         \xArray[14][18] , \xArray[14][17] , \xArray[14][16] ,
         \xArray[14][15] , \xArray[14][14] , \xArray[14][13] ,
         \xArray[14][12] , \xArray[14][11] , \xArray[14][10] , \xArray[14][9] ,
         \xArray[14][8] , \xArray[14][7] , \xArray[14][6] , \xArray[14][5] ,
         \xArray[14][4] , \xArray[14][3] , \xArray[14][2] , \xArray[14][1] ,
         \xArray[14][0] , \xArray[15][63] , \xArray[15][62] , \xArray[15][61] ,
         \xArray[15][60] , \xArray[15][59] , \xArray[15][58] ,
         \xArray[15][57] , \xArray[15][56] , \xArray[15][55] ,
         \xArray[15][54] , \xArray[15][53] , \xArray[15][52] ,
         \xArray[15][51] , \xArray[15][50] , \xArray[15][49] ,
         \xArray[15][48] , \xArray[15][47] , \xArray[15][46] ,
         \xArray[15][45] , \xArray[15][44] , \xArray[15][43] ,
         \xArray[15][42] , \xArray[15][41] , \xArray[15][40] ,
         \xArray[15][39] , \xArray[15][38] , \xArray[15][37] ,
         \xArray[15][36] , \xArray[15][35] , \xArray[15][34] ,
         \xArray[15][33] , \xArray[15][32] , \xArray[15][31] ,
         \xArray[15][30] , \xArray[15][29] , \xArray[15][28] ,
         \xArray[15][27] , \xArray[15][26] , \xArray[15][25] ,
         \xArray[15][24] , \xArray[15][23] , \xArray[15][22] ,
         \xArray[15][21] , \xArray[15][20] , \xArray[15][19] ,
         \xArray[15][18] , \xArray[15][17] , \xArray[15][16] ,
         \xArray[15][15] , \xArray[15][14] , \xArray[15][13] ,
         \xArray[15][12] , \xArray[15][11] , \xArray[15][10] , \xArray[15][9] ,
         \xArray[15][8] , \xArray[15][7] , \xArray[15][6] , \xArray[15][5] ,
         \xArray[15][4] , \xArray[15][3] , \xArray[15][2] , \xArray[15][1] ,
         \xArray[15][0] , N25537, N25538, N25539, N25540, N25541, N25542,
         N25543, N25544, N25545, N25546, N25547, N25548, N25549, N25550,
         N25551, N25552, N25553, N25554, N25555, N25556, N25557, N25558,
         N25559, N25560, N25561, N25562, N25563, N25564, N25565, N25566,
         N25567, N25568, N25569, N25570, N25571, N25572, N25573, N25574,
         N25575, N25576, N25577, N25578, N25579, N25580, N25581, N25582,
         N25583, N25584, N25601, N25602, N25603, N25604, N25605, N25606,
         N25607, N25608, N25609, N25610, N25611, N25612, N25613, N25614,
         N25615, N25616, N25617, N25618, N25619, N25620, N25621, N25622,
         N25623, N25624, N25625, N25626, N25627, N25628, N25629, N25630,
         N25631, N25632, N25633, N25634, N25635, N25636, N25637, N25638,
         N25639, N25640, N25641, N25642, N25643, N25644, N25645, N25646,
         N25647, N25648, N25649, N25650, N25651, N25652, N25653, N25654,
         N25655, N25656, N25657, N25658, N25659, N25660, N25661, N25664,
         N27809, N27810, N27811, N27812, N27813, N27814, N27815, N27816,
         N27817, N27818, N27819, N27820, N27821, N27822, N27823, N27824,
         N27825, N27826, N27827, N27828, N27829, N27830, N27831, N27832,
         N27833, N27834, N27835, N27836, N27837, N27838, N27839, N27840,
         N27841, N27842, N27843, N27844, N27845, N27846, N27847, N27848,
         N27849, N27850, N27851, N27852, N27853, N27854, N27855, N27856,
         N27857, N27858, N27859, N27860, N27861, N27862, N27863, N27864,
         N27865, N27866, N27867, N27868, N27869, N27870, N27871, N27872,
         N27873, N27874, N27875, N27876, N27877, N27878, N27879, N27880,
         N27881, N27882, N27883, N27884, N27885, N27886, N27887, N27888,
         N27889, N27890, N27891, N27892, N27893, N27894, N27895, N27896,
         N27897, N27898, N27899, N27900, N27901, N27902, N27903, N27904,
         N27905, N27906, N27907, N27908, N27909, N27910, N27911, N27912,
         N27913, N27914, N27915, N27916, N27917, N27918, N27919, N27920,
         N27921, N27922, N27923, N27924, N27925, N27926, N27927, N27928,
         N27929, N27930, N27931, N27932, N27933, N27934, N27935, N27936,
         N27937, N27938, N27939, N27940, N27941, N27942, N27943, N27944,
         N27945, N27946, N27947, N27948, N27949, N27950, N27951, N27952,
         N27953, N27954, N27955, N27956, N27957, N27958, N27959, N27960,
         N27961, N27962, N27963, N27964, N27965, N27966, N27967, N27968,
         N27969, N27970, N27971, N27972, N27973, N27974, N27975, N27976,
         N27977, N27978, N27979, N27980, N27981, N27982, N27983, N27984,
         N27985, N27986, N27987, N27988, N27989, N27990, N27991, N27992,
         N27993, N27994, N27995, N27996, N27997, N27998, N27999, N28000,
         N28001, N28002, N28003, N28004, N28005, N28006, N28007, N28008,
         N28009, N28010, N28011, N28012, N28013, N28014, N28015, N28016,
         N28017, N28018, N28019, N28020, N28021, N28022, N28023, N28024,
         N28025, N28026, N28027, N28028, N28029, N28030, N28031, N28032,
         N28033, N28034, N28035, N28036, N28037, N28038, N28039, N28040,
         N28041, N28042, N28043, N28044, N28045, N28046, N28047, N28048,
         N28049, N28050, N28051, N28052, N28053, N28054, N28055, N28056,
         N28057, N28058, N28059, N28060, N28061, N28062, N28063, N28064,
         N28065, N28066, N28067, N28068, N28069, N28070, N28071, N28072,
         N28073, N28074, N28075, N28076, N28077, N28078, N28079, N28080,
         N28081, N28082, N28083, N28084, N28085, N28086, N28087, N28088,
         N28089, N28090, N28091, N28092, N28093, N28094, N28095, N28096,
         N28097, N28098, N28099, N28100, N28101, N28102, N28103, N28104,
         N28105, N28106, N28107, N28108, N28109, N28110, N28111, N28112,
         N28113, N28114, N28115, N28116, N28117, N28118, N28119, N28120,
         N28121, N28122, N28123, N28124, N28125, N28126, N28127, N28128,
         N28129, N28130, N28131, N28132, N28133, N28134, N28135, N28136,
         N28137, N28138, N28139, N28140, N28141, N28142, N28143, N28144,
         N28145, N28146, N28147, N28148, N28149, N28150, N28151, N28152,
         N28153, N28154, N28155, N28156, N28157, N28158, N28159, N28160,
         N28161, N28162, N28163, N28164, N28165, N28166, N28167, N28168,
         N28169, N28170, N28171, N28172, N28173, N28174, N28175, N28176,
         N28177, N28178, N28179, N28180, N28181, N28182, N28183, N28184,
         N28185, N28186, N28187, N28188, N28189, N28190, N28191, N28192,
         N28193, N28194, N28195, N28196, N28197, N28198, N28199, N28200,
         N28201, N28202, N28203, N28204, N28205, N28206, N28207, N28208,
         N28209, N28210, N28211, N28212, N28213, N28214, N28215, N28216,
         N28217, N28218, N28219, N28220, N28221, N28222, N28223, N28224,
         N28225, N28226, N28227, N28228, N28229, N28230, N28231, N28232,
         N28233, N28234, N28235, N28236, N28237, N28238, N28239, N28240,
         N28241, N28242, N28243, N28244, N28245, N28246, N28247, N28248,
         N28249, N28250, N28251, N28252, N28253, N28254, N28255, N28256,
         N28257, N28258, N28259, N28260, N28261, N28262, N28263, N28264,
         N28265, N28266, N28267, N28268, N28269, N28270, N28271, N28272,
         N28273, N28274, N28275, N28276, N28277, N28278, N28279, N28280,
         N28281, N28282, N28283, N28284, N28285, N28286, N28287, N28288,
         N28289, N28290, N28291, N28292, N28293, N28294, N28295, N28296,
         N28297, N28298, N28299, N28300, N28301, N28302, N28303, N28304,
         N28305, N28306, N28307, N28308, N28309, N28310, N28311, N28312,
         N28313, N28314, N28315, N28316, N28317, N28318, N28319, N28320,
         N28321, N28322, N28323, N28324, N28325, N28326, N28327, N28328,
         N28329, N28330, N28331, N28332, N28333, N28334, N28335, N28336,
         N28337, N28338, N28339, N28340, N28341, N28342, N28343, N28344,
         N28345, N28346, N28347, N28348, N28349, N28350, N28351, N28352,
         N28353, N28354, N28355, N28356, N28357, N28358, N28359, N28360,
         N28361, N28362, N28363, N28364, N28365, N28366, N28367, N28368,
         N28369, N28370, N28371, N28372, N28373, N28374, N28375, N28376,
         N28377, N28378, N28379, N28380, N28381, N28382, N28383, N28384,
         N28385, N28386, N28387, N28388, N28389, N28390, N28391, N28392,
         N28393, N28394, N28395, N28396, N28397, N28398, N28399, N28400,
         N28401, N28402, N28403, N28404, N28405, N28406, N28407, N28408,
         N28409, N28410, N28411, N28412, N28413, N28414, N28415, N28416,
         N28417, N28418, N28419, N28420, N28421, N28422, N28423, N28424,
         N28425, N28426, N28427, N28428, N28429, N28430, N28431, N28432,
         N28433, N28434, N28435, N28436, N28437, N28438, N28439, N28440,
         N28441, N28442, N28443, N28444, N28445, N28446, N28447, N28448,
         N28449, N28450, N28451, N28452, N28453, N28454, N28455, N28456,
         N28457, N28458, N28459, N28460, N28461, N28462, N28463, N28464,
         N28465, N28466, N28467, N28468, N28469, N28470, N28471, N28472,
         N28473, N28474, N28475, N28476, N28477, N28478, N28479, N28480,
         N28481, N28482, N28483, N28484, N28485, N28486, N28487, N28488,
         N28489, N28490, N28491, N28492, N28493, N28494, N28495, N28496,
         N28497, N28498, N28499, N28500, N28501, N28502, N28503, N28504,
         N28505, N28506, N28507, N28508, N28509, N28510, N28511, N28512,
         N28513, N28514, N28515, N28516, N28517, N28518, N28519, N28520,
         N28521, N28522, N28523, N28524, N28525, N28526, N28527, N28528,
         N28529, N28530, N28531, N28532, N28533, N28534, N28535, N28536,
         N28537, N28538, N28539, N28540, N28541, N28542, N28543, N28544,
         N28545, N28546, N28547, N28548, N28549, N28550, N28551, N28552,
         N28553, N28554, N28555, N28556, N28557, N28558, N28559, N28560,
         N28561, N28562, N28563, N28564, N28565, N28566, N28567, N28568,
         N28569, N28570, N28571, N28572, N28573, N28574, N28575, N28576,
         N28577, N28578, N28579, N28580, N28581, N28582, N28583, N28584,
         N28585, N28586, N28587, N28588, N28589, N28590, N28591, N28592,
         N28593, N28594, N28595, N28596, N28597, N28598, N28599, N28600,
         N28601, N28602, N28603, N28604, N28605, N28606, N28607, N28608,
         N28609, N28610, N28611, N28612, N28613, N28614, N28615, N28616,
         N28617, N28618, N28619, N28620, N28621, N28622, N28623, N28624,
         N28625, N28626, N28627, N28628, N28629, N28630, N28631, N28632,
         N28633, N28634, N28635, N28636, N28637, N28638, N28639, N28640,
         N28641, N28642, N28643, N28644, N28645, N28646, N28647, N28648,
         N28649, N28650, N28651, N28652, N28653, N28654, N28655, N28656,
         N28657, N28658, N28659, N28660, N28661, N28662, N28663, N28664,
         N28665, N28666, N28667, N28668, N28669, N28670, N28671, N28672,
         N28673, N28674, N28675, N28676, N28677, N28678, N28679, N28680,
         N28681, N28682, N28683, N28684, N28685, N28686, N28687, N28688,
         N28689, N28690, N28691, N28692, N28693, N28694, N28695, N28696,
         N28697, N28698, N28699, N28700, N28701, N28702, N28703, N28704,
         N28705, N28706, N28707, N28708, N28709, N28710, N28711, N28712,
         N28713, N28714, N28715, N28716, N28717, N28718, N28719, N28720,
         N28721, N28722, N28723, N28724, N28725, N28726, N28727, N28728,
         N28729, N28730, N28731, N28732, N28733, N28734, N28735, N28736,
         N28737, N28738, N28739, N28740, N28741, N28742, N28743, N28744,
         N28745, N28746, N28747, N28748, N28749, N28750, N28751, N28752,
         N28753, N28754, N28755, N28756, N28757, N28758, N28759, N28760,
         N28761, N28762, N28763, N28764, N28765, N28766, N28767, N28768,
         N28769, N28770, N28771, N28772, N28773, N28774, N28775, N28776,
         N28777, N28778, N28779, N28780, N28781, N28782, N28783, N28784,
         N28785, N28786, N28787, N28788, N28789, N28790, N28791, N28792,
         N28793, N28794, N28795, N28796, N28797, N28798, N28799, N28800,
         N28801, N28802, N28803, N28804, N28805, N28806, N28807, N28808,
         N28809, N28810, N28811, N28812, N28813, N28814, N28815, N28816,
         N28817, N28818, N28819, N28820, N28821, N28822, N28823, N28824,
         N28825, N28826, N28827, N28828, N28829, N28830, N28831, N28832,
         N28833, N28834, N28835, N28836, N28837, N28838, N28839, N28840,
         N28841, N28842, N28843, N28844, N28845, N28846, N28847, N28848,
         N28849, N28850, N28851, N28852, N28853, N28854, N28855, N28856,
         N28857, N28858, N28859, N28860, N28861, N28862, N28863, N28864,
         N28865, N28866, N28867, N28868, N28869, N28870, N28871, N28872,
         N28873, N28874, N28875, N28876, N28877, N28878, N28879, N28880,
         N29546, N29547, N29548, N29549, N29550, N29551, N29552, N29553,
         N29554, N29555, N29556, N29557, N29558, N29559, N29560, N29561,
         N29562, N29563, N29564, N29565, N29566, N29567, N29568, N29569,
         N29570, N29571, N29572, N29573, N29574, N29575, N29576, N29577,
         N29578, N29579, N29580, N29581, N29582, N29583, N29584, N29585,
         N29586, N29587, N29588, N29589, N29590, N29591, N29592, N29593,
         N29594, N29595, N29596, N29597, N29598, N29599, N29600, N29601,
         N29602, N29603, N29604, N29605, N29606, N29607, N29608, N29609,
         N29610, N29611, N29612, N29613, N29614, N29615, N29616, N29617,
         N29618, N29619, N29620, N29621, N29622, N29623, N29624, N29625,
         N29626, N29627, N29628, N29629, N29630, N29631, N29632, N29633,
         N29634, N29635, N29636, N29637, N29638, N29639, N29640, N29641,
         N29642, N29643, N29644, N29645, N29646, N29647, N29648, N29649,
         N29650, N29651, N29652, N29653, N29654, N29655, N29656, N29657,
         N29658, N29659, N29660, N29661, N29662, N29663, N29664, N29665,
         N29666, N29667, N29668, N29669, N29670, N29671, N29672, N29673,
         N30314, N30315, N30316, N30317, N30318, N30319, N30320, N30321,
         N30322, N30323, N30324, N30325, N30326, N30327, N30328, N30329,
         N30330, N30331, N30332, N30333, N30334, N30335, N30336, N30337,
         N30338, N30339, N30340, N30341, N30342, N30343, N30344, N30345,
         N30346, N30347, N30348, N30349, N30350, N30351, N30352, N30353,
         N30354, N30355, N30356, N30357, N30358, N30359, N30360, N30361,
         N30362, N30363, N30364, N30365, N30366, N30367, N30368, N30369,
         N30370, N30371, N30372, N30373, N30374, N30375, N30376, N30377,
         N30378, N30379, N30380, N30381, N30382, N30383, N30384, N30385,
         N30386, N30387, N30388, N30389, N30390, N30391, N30392, N30393,
         N30394, N30395, N30396, N30397, N30398, N30399, N30400, N30401,
         N30402, N30403, N30404, N30405, N30406, N30407, N30408, N30409,
         N30410, N30411, N30412, N30413, N30414, N30415, N30416, N30417,
         N30418, N30419, N30420, N30421, N30422, N30423, N30424, N30425,
         N30426, N30427, N30428, N30429, N30430, N30431, N30432, N30433,
         N30434, N30435, N30436, N30437, N30438, N30439, N30440, N30441,
         N31274, N31275, N31276, N31277, N31278, N31279, N31280, N31281,
         N31282, N31283, N31284, N31285, N31286, N31287, N31288, N31289,
         N31290, N31291, N31292, N31293, N31294, N31295, N31296, N31297,
         N31298, N31299, N31300, N31301, N31302, N31303, N31304, N31305,
         N31306, N31307, N31308, N31309, N31310, N31311, N31312, N31313,
         N31314, N31315, N31316, N31317, N31318, N31319, N31320, N31321,
         N31322, N31323, N31324, N31325, N31326, N31327, N31328, N31329,
         N31330, N31331, N31332, N31333, N31334, N31335, N31336, N31337,
         N31338, N31339, N31340, N31341, N31342, N31343, N31344, N31345,
         N31346, N31347, N31348, N31349, N31350, N31351, N31352, N31353,
         N31354, N31355, N31356, N31357, N31358, N31359, N31360, N31361,
         N31362, N31363, N31364, N31365, N31366, N31367, N31368, N31369,
         N31370, N31371, N31372, N31373, N31374, N31375, N31376, N31377,
         N31378, N31379, N31380, N31381, N31382, N31383, N31384, N31385,
         N31386, N31387, N31388, N31389, N31390, N31391, N31392, N31393,
         N31394, N31395, N31396, N31397, N31398, N31399, N31400, N31401,
         N31850, N31851, N31852, N31853, N31854, N31855, N31856, N31857,
         N31858, N31859, N31860, N31861, N31862, N31863, N31864, N31865,
         N31866, N31867, N31868, N31869, N31870, N31871, N31872, N31873,
         N31874, N31875, N31876, N31877, N31878, N31879, N31880, N31881,
         N31882, N31883, N31884, N31885, N31886, N31887, N31888, N31889,
         N31890, N31891, N31892, N31893, N31894, N31895, N31896, N31897,
         N31898, N31899, N31900, N31901, N31902, N31903, N31904, N31905,
         N31906, N31907, N31908, N31909, N31910, N31911, N31912, N31913,
         N31914, N31915, N31916, N31917, N31918, N31919, N31920, N31921,
         N31922, N31923, N31924, N31925, N31926, N31927, N31928, N31929,
         N31930, N31931, N31932, N31933, N31934, N31935, N31936, N31937,
         N31938, N31939, N31940, N31941, N31942, N31943, N31944, N31945,
         N31946, N31947, N31948, N31949, N31950, N31951, N31952, N31953,
         N31954, N31955, N31956, N31957, N31958, N31959, N31960, N31961,
         N31962, N31963, N31964, N31965, N31966, N31967, N31968, N31969,
         N31970, N31971, N31972, N31973, N31974, N31975, N31976, N31977,
         N32618, N32619, N32620, N32621, N32622, N32623, N32624, N32625,
         N32626, N32627, N32628, N32629, N32630, N32631, N32632, N32633,
         N32634, N32635, N32636, N32637, N32638, N32639, N32640, N32641,
         N32642, N32643, N32644, N32645, N32646, N32647, N32648, N32649,
         N32650, N32651, N32652, N32653, N32654, N32655, N32656, N32657,
         N32658, N32659, N32660, N32661, N32662, N32663, N32664, N32665,
         N32666, N32667, N32668, N32669, N32670, N32671, N32672, N32673,
         N32674, N32675, N32676, N32677, N32678, N32679, N32680, N32681,
         N32682, N32683, N32684, N32685, N32686, N32687, N32688, N32689,
         N32690, N32691, N32692, N32693, N32694, N32695, N32696, N32697,
         N32698, N32699, N32700, N32701, N32702, N32703, N32704, N32705,
         N32706, N32707, N32708, N32709, N32710, N32711, N32712, N32713,
         N32714, N32715, N32716, N32717, N32718, N32719, N32720, N32721,
         N32722, N32723, N32724, N32725, N32726, N32727, N32728, N32729,
         N32730, N32731, N32732, N32733, N32734, N32735, N32736, N32737,
         N32738, N32739, N32740, N32741, N32742, N32743, N32744, N32745,
         N33578, N33579, N33580, N33581, N33582, N33583, N33584, N33585,
         N33586, N33587, N33588, N33589, N33590, N33591, N33592, N33593,
         N33594, N33595, N33596, N33597, N33598, N33599, N33600, N33601,
         N33602, N33603, N33604, N33605, N33606, N33607, N33608, N33609,
         N33610, N33611, N33612, N33613, N33614, N33615, N33616, N33617,
         N33618, N33619, N33620, N33621, N33622, N33623, N33624, N33625,
         N33626, N33627, N33628, N33629, N33630, N33631, N33632, N33633,
         N33634, N33635, N33636, N33637, N33638, N33639, N33640, N33641,
         N33642, N33643, N33644, N33645, N33646, N33647, N33648, N33649,
         N33650, N33651, N33652, N33653, N33654, N33655, N33656, N33657,
         N33658, N33659, N33660, N33661, N33662, N33663, N33664, N33665,
         N33666, N33667, N33668, N33669, N33670, N33671, N33672, N33673,
         N33674, N33675, N33676, N33677, N33678, N33679, N33680, N33681,
         N33682, N33683, N33684, N33685, N33686, N33687, N33688, N33689,
         N33690, N33691, N33692, N33693, N33694, N33695, N33696, N33697,
         N33698, N33699, N33700, N33701, N33702, N33703, N33704, N33705,
         N33706, N33707, N33708, N33709, N33710, N33711, N33712, N33713,
         N33714, N33715, N33716, N33717, N33718, N33719, N33720, N33721,
         N33722, N33723, N33724, N33725, N33726, N33727, N33728, N33729,
         N33730, N33731, N33732, N33733, N33734, N33735, N33736, N33737,
         N33738, N33739, N33740, N33741, N33742, N33743, N33744, N33745,
         N33746, N33747, N33748, N33749, N33750, N33751, N33752, N33753,
         N33754, N33755, N33756, N33757, N33758, N33759, N33760, N33761,
         N33762, N33763, N33764, N33765, N33766, N33767, N33768, N33769,
         N33770, N33771, N33772, N33773, N33774, N33775, N33776, N33777,
         N33778, N33779, N33780, N33781, N33782, N33783, N33784, N33785,
         N33786, N33787, N33788, N33789, N33790, N33791, N33792, N33793,
         N33794, N33795, N33796, N33797, N33798, N33799, N33800, N33801,
         N33802, N33803, N33804, N33805, N33806, N33807, N33808, N33809,
         N33810, N33811, N33812, N33813, N33814, N33815, N33816, N33817,
         N33818, N33819, N33820, N33821, N33822, N33823, N33824, N33825,
         N33826, N33827, N33828, N33829, N33830, N33831, N33832, N33833,
         N33834, N33835, N33836, N33837, N33838, N33839, N33840, N33841,
         N33842, N33843, N33844, N33845, N33846, N33847, N33848, N33849,
         N33850, N33851, N33852, N33853, N33854, N33855, N33856, N33857,
         N33858, N33859, N33860, N33861, N33862, N33863, N33864, N33865,
         N33866, N33867, N33868, N33869, N33870, N33871, N33872, N33873,
         N33874, N33875, N33876, N33877, N33878, N33879, N33880, N33881,
         N33882, N33883, N33884, N33885, N33886, N33887, N33888, N33889,
         N33890, N33891, N33892, N33893, N33894, N33895, N33896, N33897,
         N33898, N33899, N33900, N33901, N33902, N33903, N33904, N33905,
         N33906, N33907, N33908, N33909, N33910, N33911, N33912, N33913,
         N33914, N33915, N33916, N33917, N33918, N33919, N33920, N33921,
         N33922, N33923, N33924, N33925, N33926, N33927, N33928, N33929,
         N33930, N33931, N33932, N33933, N33934, N33935, N33936, N33937,
         N33938, N33939, N33940, N33941, N33942, N33943, N33944, N33945,
         N33946, N33947, N33948, N33949, N33950, N33951, N33952, N33953,
         N33954, N33955, N33956, N33957, N33958, N33959, N33960, N33961,
         N33962, N33963, N33964, N33965, N33966, N33967, N33968, N33969,
         N33970, N33971, N33972, N33973, N33974, N33975, N33976, N33977,
         N33978, N33979, N33980, N33981, N33982, N33983, N33984, N33985,
         N33986, N33987, N33988, N33989, N33990, N33991, N33992, N33993,
         N33994, N33995, N33996, N33997, N33998, N33999, N34000, N34001,
         N34002, N34003, N34004, N34005, N34006, N34007, N34008, N34009,
         N34010, N34011, N34012, N34013, N34014, N34015, N34016, N34017,
         N34018, N34019, N34020, N34021, N34022, N34023, N34024, N34025,
         N34026, N34027, N34028, N34029, N34030, N34031, N34032, N34033,
         N34034, N34035, N34036, N34037, N34038, N34039, N34040, N34041,
         N34042, N34043, N34044, N34045, N34046, N34047, N34048, N34049,
         N34050, N34051, N34052, N34053, N34054, N34055, N34056, N34057,
         N34058, N34059, N34060, N34061, N34062, N34063, N34064, N34065,
         N34066, N34067, N34068, N34069, N34070, N34071, N34072, N34073,
         N34074, N34075, N34076, N34077, N34078, N34079, N34080, N34081,
         N34082, N34083, N34084, N34085, N34086, N34087, N34088, N34089,
         N34666, N34667, N34668, N34669, N34670, N34671, N34672, N34673,
         N34674, N34675, N34676, N34677, N34678, N34679, N34680, N34681,
         N34682, N34683, N34684, N34685, N34686, N34687, N34688, N34689,
         N34690, N34691, N34692, N34693, N34694, N34695, N34696, N34697,
         N34698, N34699, N34700, N34701, N34702, N34703, N34704, N34705,
         N34706, N34707, N34708, N34709, N34710, N34711, N34712, N34713,
         N34714, N34715, N34716, N34717, N34718, N34719, N34720, N34721,
         N34722, N34723, N34724, N34725, N34726, N34727, N34728, N34729,
         N34730, N34731, N34732, N34733, N34734, N34735, N34736, N34737,
         N34738, N34739, N34740, N34741, N34742, N34743, N34744, N34745,
         N34746, N34747, N34748, N34749, N34750, N34751, N34752, N34753,
         N34754, N34755, N34756, N34757, N34758, N34759, N34760, N34761,
         N34762, N34763, N34764, N34765, N34766, N34767, N34768, N34769,
         N34770, N34771, N34772, N34773, N34774, N34775, N34776, N34777,
         N34778, N34779, N34780, N34781, N34782, N34783, N34784, N34785,
         N34786, N34787, N34788, N34789, N34790, N34791, N34792, N34793,
         N34877, N34878, N34879, N34880, N34881, N34882, N34883, N34884,
         N34885, N34886, N34887, N34888, N34889, N34890, N34891, N34892,
         N34893, N34894, N34895, N34896, N34897, N34898, N34899, N34900,
         N34901, N34902, N34903, N34904, N34905, N34906, N34907, N34908,
         N34910, N34911, N34912, N34913, N34914, N34915, N34916, N34917,
         N34918, N34919, N34920, N34921, N34922, N34923, N34924, N34925,
         N34926, N34927, N34928, N34929, N34930, N34931, N34932, N34933,
         N34934, N34935, N34936, N34937, N34938, N34939, N34940, N34941,
         N34942, N34943, N34944, N34945, N34946, N34947, N34948, N34949,
         N34950, N34951, N34952, N34953, N34954, N34955, N34956, N34957,
         N34958, N34959, N34960, N34961, N34962, N34963, N34964, N34965,
         N34966, N34967, N34968, N34969, N34970, N34971, N34972, N34973,
         N34983, N35017, N35018, N35019, N35020, N35021, N35022, N35023,
         N35024, N35025, N35026, N35027, N35028, N35029, N35030, N35031,
         N35032, N35033, N35034, N35035, N35036, N35037, N35038, N35039,
         N35040, N35041, N35042, N35043, N35044, N35045, N35046, N35047,
         N35048, N35084, N35085, N35086, N35087, N35088, N35089, N35090,
         N35091, N35092, N35093, N35094, N35095, N35096, N35097, N35098,
         N35099, N35100, N35101, N35102, N35103, N35104, N35105, N35106,
         N35107, N35108, N35109, N35110, N35111, N35112, N35113, N35114,
         N35115, N35189, N35192, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n109,
         n110, n111, n112, n116, n117, n118, n119, n123, n124, n125, n126,
         n130, n131, n132, n133, n135, n159, n160, n161, n164, n165, n181,
         n183, n184, n185, n187, n188, n189, n191, n192, n193, n195, n196,
         n197, n199, n200, n201, n203, n204, n205, n207, n208, n209, n211,
         n212, n213, n215, n216, n218, n219, n220, n222, n223, n224, n226,
         n227, n228, n230, n231, n232, n234, n235, n236, n238, n239, n240,
         n241, n242, n243, n244, n248, n249, n250, n251, n252, n253, n254,
         n255, n257, n258, n261, n262, n266, n267, n268, n269, n271, n272,
         n273, n274, n277, n278, n279, n280, n281, n282, n285, n286, n287,
         n288, n289, n290, n293, n294, n295, n296, n297, n298, n301, n302,
         n303, n304, n305, n306, n309, n310, n311, n312, n313, n314, n317,
         n318, n319, n320, n321, n322, n325, n326, n327, n328, n329, n330,
         n333, n334, n335, n336, n337, n338, n341, n342, n343, n344, n345,
         n346, n349, n350, n351, n352, n353, n354, n357, n358, n359, n360,
         n361, n362, n365, n366, n367, n368, n369, n370, n373, n374, n375,
         n376, n377, n378, n381, n382, n383, n384, n385, n386, n389, n390,
         n391, n392, n393, n394, n397, n398, n399, n400, n401, n402, n405,
         n406, n407, n408, n409, n410, n413, n414, n415, n416, n417, n418,
         n421, n422, n423, n424, n425, n426, n429, n430, n431, n432, n433,
         n434, n437, n438, n439, n440, n441, n442, n445, n446, n447, n448,
         n449, n450, n453, n454, n455, n456, n457, n458, n461, n462, n463,
         n464, n465, n466, n469, n470, n471, n472, n473, n474, n477, n478,
         n479, n480, n481, n482, n485, n486, n487, n488, n489, n490, n493,
         n494, n495, n496, n497, n498, n501, n502, n503, n504, n505, n506,
         n509, n510, n511, n512, n513, n514, n517, n518, n519, n520, n521,
         n522, n525, n526, n527, n528, n529, n530, n533, n534, n535, n536,
         n537, n538, n541, n542, n543, n544, n545, n546, n549, n550, n551,
         n552, n553, n554, n557, n558, n559, n560, n561, n562, n565, n566,
         n567, n568, n569, n570, n573, n574, n575, n576, n577, n578, n581,
         n582, n583, n584, n585, n586, n589, n590, n591, n592, n593, n594,
         n597, n598, n599, n600, n601, n602, n605, n606, n607, n608, n609,
         n610, n613, n614, n615, n616, n617, n618, n621, n622, n623, n624,
         n625, n626, n629, n630, n631, n632, n633, n634, n637, n638, n639,
         n640, n641, n642, n645, n646, n647, n648, n649, n650, n653, n654,
         n655, n656, n657, n658, n661, n662, n663, n664, n665, n666, n669,
         n670, n671, n672, n673, n674, n677, n678, n679, n680, n681, n682,
         n685, n686, n687, n688, n689, n690, n693, n694, n695, n696, n697,
         n698, n701, n702, n703, n704, n705, n706, n709, n710, n711, n712,
         n713, n714, n717, n718, n719, n720, n721, n722, n725, n726, n727,
         n728, n729, n730, n733, n734, n735, n736, n737, n738, n741, n742,
         n743, n744, n745, n746, n749, n750, n751, n752, n753, n754, n757,
         n758, n759, n760, n761, n762, n765, n766, n767, n768, n769, n770,
         n773, n775, n777, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n981, n982, n983, n984, n986,
         n987, n988, n989, n991, n992, n993, n994, n996, n997, n998, n999,
         n1001, n1002, n1003, n1004, n1006, n1007, n1008, n1009, n1011, n1012,
         n1013, n1014, n1016, n1017, n1018, n1019, n1021, n1022, n1023, n1024,
         n1026, n1027, n1028, n1029, n1031, n1032, n1033, n1034, n1036, n1037,
         n1038, n1039, n1041, n1042, n1043, n1044, n1046, n1047, n1048, n1049,
         n1051, n1052, n1053, n1054, n1056, n1057, n1058, n1059, n1061, n1062,
         n1063, n1064, n1066, n1067, n1068, n1069, n1071, n1072, n1073, n1074,
         n1076, n1077, n1078, n1079, n1081, n1082, n1083, n1084, n1086, n1087,
         n1088, n1089, n1091, n1092, n1093, n1094, n1096, n1097, n1098, n1099,
         n1101, n1102, n1103, n1104, n1106, n1107, n1108, n1109, n1111, n1112,
         n1113, n1114, n1116, n1117, n1118, n1119, n1121, n1122, n1123, n1124,
         n1126, n1127, n1128, n1129, n1131, n1132, n1133, n1134, n1136, n1137,
         n1138, n1139, n1141, n1142, n1143, n1144, n1146, n1147, n1148, n1149,
         n1151, n1152, n1153, n1154, n1156, n1157, n1158, n1159, n1161, n1162,
         n1163, n1164, n1166, n1167, n1168, n1169, n1171, n1172, n1173, n1174,
         n1176, n1177, n1178, n1179, n1181, n1182, n1183, n1184, n1186, n1187,
         n1188, n1189, n1191, n1192, n1193, n1194, n1196, n1197, n1198, n1199,
         n1201, n1202, n1203, n1204, n1206, n1207, n1208, n1209, n1211, n1212,
         n1213, n1214, n1216, n1217, n1218, n1219, n1221, n1222, n1223, n1224,
         n1226, n1227, n1228, n1229, n1231, n1232, n1233, n1234, n1236, n1237,
         n1238, n1239, n1241, n1242, n1243, n1244, n1246, n1247, n1248, n1249,
         n1251, n1252, n1253, n1254, n1256, n1257, n1258, n1259, n1261, n1262,
         n1263, n1264, n1266, n1267, n1268, n1269, n1271, n1272, n1273, n1274,
         n1276, n1277, n1278, n1279, n1281, n1282, n1283, n1284, n1286, n1287,
         n1288, n1289, n1292, n1293, n1294, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1751, n1753,
         n1755, n1756, n1757, n1758, n1759, n1762, n1764, n1765, n1766, n1767,
         n1768, n1771, n1773, n1774, n1775, n1776, n1777, n1780, n1782, n1783,
         n1784, n1785, n1786, n1789, n1791, n1792, n1793, n1794, n1795, n1798,
         n1800, n1801, n1802, n1803, n1804, n1807, n1809, n1810, n1811, n1812,
         n1813, n1816, n1818, n1819, n1820, n1821, n1822, n1825, n1827, n1828,
         n1829, n1830, n1831, n1834, n1836, n1837, n1838, n1839, n1840, n1843,
         n1845, n1846, n1847, n1848, n1849, n1852, n1854, n1855, n1856, n1857,
         n1858, n1861, n1863, n1864, n1865, n1866, n1867, n1870, n1872, n1873,
         n1874, n1875, n1876, n1879, n1881, n1882, n1883, n1884, n1885, n1888,
         n1890, n1891, n1892, n1893, n1894, n1897, n1899, n1900, n1901, n1902,
         n1903, n1906, n1908, n1909, n1910, n1911, n1912, n1915, n1917, n1918,
         n1919, n1920, n1921, n1924, n1926, n1927, n1928, n1929, n1930, n1933,
         n1935, n1936, n1937, n1938, n1939, n1942, n1944, n1945, n1946, n1947,
         n1948, n1951, n1953, n1954, n1955, n1956, n1957, n1960, n1962, n1963,
         n1964, n1965, n1966, n1969, n1971, n1972, n1973, n1974, n1975, n1978,
         n1980, n1981, n1982, n1983, n1984, n1987, n1989, n1990, n1991, n1992,
         n1993, n1996, n1998, n1999, n2000, n2001, n2002, n2005, n2007, n2008,
         n2009, n2010, n2011, n2014, n2016, n2017, n2018, n2019, n2020, n2023,
         n2025, n2026, n2027, n2028, n2029, n2032, n2034, n2035, n2036, n2037,
         n2038, n2041, n2043, n2044, n2045, n2046, n2047, n2050, n2052, n2053,
         n2054, n2055, n2056, n2059, n2061, n2062, n2063, n2064, n2065, n2068,
         n2070, n2071, n2072, n2073, n2074, n2077, n2079, n2080, n2081, n2082,
         n2083, n2086, n2088, n2089, n2090, n2091, n2092, n2095, n2097, n2098,
         n2099, n2100, n2101, n2104, n2106, n2107, n2108, n2109, n2110, n2113,
         n2115, n2116, n2117, n2118, n2119, n2122, n2124, n2125, n2126, n2127,
         n2128, n2131, n2133, n2134, n2135, n2136, n2137, n2140, n2142, n2143,
         n2144, n2145, n2146, n2149, n2151, n2152, n2153, n2154, n2155, n2158,
         n2160, n2161, n2162, n2163, n2164, n2167, n2169, n2170, n2171, n2172,
         n2173, n2176, n2178, n2179, n2180, n2181, n2182, n2185, n2187, n2188,
         n2189, n2190, n2191, n2194, n2196, n2197, n2198, n2199, n2200, n2203,
         n2205, n2206, n2207, n2208, n2209, n2212, n2214, n2215, n2216, n2217,
         n2218, n2221, n2223, n2224, n2225, n2226, n2227, n2230, n2232, n2233,
         n2234, n2235, n2236, n2239, n2241, n2242, n2243, n2244, n2245, n2248,
         n2250, n2251, n2252, n2253, n2254, n2257, n2259, n2260, n2261, n2262,
         n2263, n2266, n2268, n2269, n2270, n2271, n2272, n2275, n2277, n2278,
         n2279, n2280, n2281, n2284, n2286, n2287, n2288, n2289, n2290, n2293,
         n2295, n2296, n2297, n2298, n2299, n2302, n2304, n2305, n2306, n2307,
         n2308, n2311, n2313, n2314, n2315, n2316, n2317, n2323, n2325, n2326,
         n2327, n2328, n2331, n2334, n2335, n2337, n2338, n2340, n2341, n2343,
         n2344, n2346, n2347, n2349, n2350, n2352, n2353, n2355, n2356, n2358,
         n2359, n2361, n2362, n2364, n2365, n2367, n2368, n2370, n2371, n2373,
         n2374, n2376, n2377, n2379, n2380, n2382, n2383, n2385, n2386, n2388,
         n2389, n2392, n2394, n2395, n2397, n2398, n2400, n2401, n2403, n2404,
         n2406, n2407, n2409, n2410, n2412, n2413, n2415, n2416, n2418, n2419,
         n2421, n2422, n2424, n2425, n2427, n2428, n2430, n2431, n2433, n2434,
         n2436, n2437, n2439, n2440, n2442, n2443, n2445, n2446, n2448, n2449,
         n2451, n2452, n2454, n2455, n2457, n2458, n2460, n2461, n2463, n2464,
         n2466, n2467, n2469, n2470, n2472, n2473, n2475, n2476, n2478, n2479,
         n2481, n2482, n2484, n2485, n2487, n2488, n2490, n2491, n2493, n2494,
         n2496, n2497, n2499, n2500, n2502, n2503, n2505, n2506, n2508, n2509,
         n2511, n2512, n2514, n2515, n2517, n2518, n2520, n2521, n2523, n2524,
         n2526, n2528, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2805,
         n2806, n2808, n2809, n2811, n2813, n2815, n2817, n2819, n2821, n2823,
         n2825, n2827, n2829, n2831, n2833, n2835, n2837, n2839, n2841, n2843,
         n2845, n2847, n2849, n2851, n2853, n2855, n2857, n2859, n2861, n2863,
         n2865, n2867, n2869, n2871, n2873, n2875, n2877, n2879, n2881, n2883,
         n2885, n2887, n2889, n2891, n2893, n2895, n2897, n2899, n2901, n2903,
         n2905, n2907, n2909, n2911, n2913, n2915, n2917, n2919, n2921, n2923,
         n2925, n2927, n2929, n2931, n2933, n2935, n2936, n2937, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3010, n3011, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3080, n3081, n3082, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3295, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3362, n3363, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3431, n3432, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3500, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3651, n3652, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3665, n3667, n3668, n3669, n3671, n3674, n3675, n3676,
         n3678, n3680, n3682, n3685, n3687, n3689, n3691, n3693, n3695, n3696,
         n3697, n3699, n3700, n3703, n3705, n3706, n3707, n3708, n3709, n3711,
         n3714, n3717, n3718, n3719, n3720, n3721, n3723, n3724, n3725, n3726,
         n3727, n3729, n3732, n3735, n3736, n3737, n3738, n3739, n3741, n3742,
         n3743, n3744, n3745, n3747, n3750, n3753, n3754, n3755, n3756, n3757,
         n3759, n3760, n3761, n3762, n3763, n3765, n3768, n3771, n3772, n3773,
         n3774, n3775, n3777, n3778, n3779, n3780, n3781, n3783, n3786, n3789,
         n3790, n3791, n3792, n3793, n3795, n3796, n3797, n3798, n3799, n3801,
         n3804, n3807, n3808, n3809, n3810, n3811, n3813, n3814, n3815, n3816,
         n3817, n3819, n3822, n3825, n3826, n3827, n3828, n3829, n3831, n3832,
         n3833, n3834, n3835, n3837, n3840, n3843, n3844, n3845, n3846, n3847,
         n3849, n3850, n3851, n3852, n3853, n3855, n3858, n3861, n3862, n3863,
         n3864, n3865, n3867, n3868, n3869, n3870, n3871, n3873, n3876, n3879,
         n3880, n3881, n3882, n3883, n3885, n3886, n3887, n3888, n3889, n3891,
         n3894, n3897, n3898, n3899, n3900, n3901, n3903, n3904, n3905, n3906,
         n3907, n3909, n3912, n3915, n3916, n3917, n3918, n3919, n3921, n3922,
         n3923, n3924, n3925, n3927, n3930, n3933, n3934, n3935, n3936, n3937,
         n3939, n3940, n3941, n3942, n3943, n3945, n3948, n3951, n3952, n3953,
         n3954, n3955, n3957, n3958, n3959, n3960, n3961, n3963, n3966, n3969,
         n3970, n3971, n3972, n3973, n3975, n3976, n3977, n3978, n3979, n3981,
         n3984, n3987, n3988, n3989, n3990, n3991, n3993, n3994, n3995, n3996,
         n3997, n3999, n4002, n4005, n4006, n4007, n4008, n4009, n4011, n4012,
         n4013, n4014, n4015, n4017, n4020, n4023, n4024, n4025, n4026, n4027,
         n4029, n4030, n4031, n4032, n4033, n4035, n4038, n4041, n4042, n4043,
         n4044, n4045, n4047, n4048, n4049, n4050, n4051, n4053, n4056, n4059,
         n4060, n4061, n4062, n4063, n4065, n4066, n4067, n4068, n4069, n4071,
         n4074, n4077, n4078, n4079, n4080, n4081, n4083, n4084, n4085, n4086,
         n4087, n4089, n4092, n4095, n4096, n4097, n4098, n4099, n4101, n4102,
         n4103, n4104, n4105, n4107, n4110, n4113, n4114, n4115, n4116, n4117,
         n4119, n4120, n4121, n4122, n4123, n4125, n4128, n4131, n4132, n4133,
         n4134, n4135, n4137, n4138, n4139, n4140, n4141, n4143, n4146, n4149,
         n4150, n4151, n4152, n4153, n4155, n4156, n4157, n4158, n4159, n4161,
         n4164, n4167, n4168, n4169, n4170, n4171, n4173, n4174, n4175, n4176,
         n4177, n4179, n4182, n4185, n4186, n4187, n4188, n4189, n4191, n4192,
         n4193, n4194, n4195, n4197, n4200, n4203, n4204, n4205, n4206, n4207,
         n4209, n4210, n4211, n4212, n4213, n4215, n4218, n4221, n4222, n4223,
         n4224, n4225, n4227, n4228, n4229, n4230, n4231, n4233, n4236, n4239,
         n4240, n4241, n4242, n4243, n4245, n4246, n4247, n4248, n4249, n4251,
         n4254, n4257, n4258, n4259, n4260, n4261, n4263, n4264, n4265, n4266,
         n4267, n4269, n4272, n4275, n4276, n4277, n4278, n4279, n4281, n4282,
         n4283, n4284, n4285, n4287, n4290, n4293, n4294, n4295, n4296, n4297,
         n4299, n4300, n4301, n4302, n4303, n4305, n4308, n4311, n4312, n4313,
         n4314, n4315, n4317, n4318, n4319, n4320, n4321, n4323, n4326, n4329,
         n4330, n4331, n4332, n4333, n4335, n4336, n4337, n4338, n4339, n4341,
         n4344, n4347, n4348, n4349, n4350, n4351, n4353, n4354, n4355, n4356,
         n4357, n4359, n4362, n4365, n4366, n4367, n4368, n4369, n4371, n4372,
         n4373, n4374, n4375, n4377, n4380, n4383, n4384, n4385, n4386, n4387,
         n4389, n4390, n4391, n4392, n4393, n4395, n4398, n4401, n4402, n4403,
         n4404, n4405, n4407, n4408, n4409, n4410, n4411, n4413, n4416, n4419,
         n4420, n4421, n4422, n4423, n4425, n4426, n4427, n4428, n4429, n4431,
         n4434, n4437, n4438, n4439, n4440, n4441, n4443, n4444, n4445, n4446,
         n4447, n4449, n4452, n4455, n4456, n4457, n4458, n4459, n4461, n4462,
         n4463, n4464, n4465, n4467, n4470, n4473, n4474, n4475, n4476, n4477,
         n4479, n4480, n4481, n4482, n4483, n4485, n4488, n4491, n4492, n4493,
         n4494, n4495, n4497, n4498, n4499, n4500, n4501, n4503, n4506, n4509,
         n4510, n4511, n4512, n4513, n4515, n4516, n4517, n4518, n4519, n4521,
         n4524, n4527, n4528, n4529, n4530, n4531, n4533, n4534, n4535, n4536,
         n4537, n4539, n4542, n4545, n4546, n4547, n4548, n4549, n4551, n4552,
         n4553, n4554, n4555, n4557, n4560, n4563, n4564, n4565, n4566, n4567,
         n4569, n4570, n4571, n4572, n4573, n4575, n4578, n4581, n4582, n4583,
         n4584, n4585, n4587, n4588, n4589, n4590, n4591, n4593, n4596, n4599,
         n4600, n4601, n4602, n4603, n4605, n4606, n4607, n4608, n4609, n4611,
         n4614, n4617, n4618, n4619, n4620, n4621, n4623, n4624, n4625, n4626,
         n4627, n4629, n4632, n4635, n4636, n4637, n4638, n4639, n4641, n4642,
         n4643, n4644, n4645, n4647, n4650, n4653, n4654, n4655, n4656, n4657,
         n4659, n4660, n4661, n4662, n4663, n4665, n4668, n4671, n4672, n4673,
         n4674, n4675, n4677, n4678, n4679, n4680, n4681, n4683, n4686, n4689,
         n4690, n4691, n4692, n4693, n4695, n4696, n4697, n4698, n4699, n4701,
         n4704, n4707, n4708, n4709, n4710, n4711, n4713, n4714, n4715, n4716,
         n4717, n4719, n4722, n4725, n4726, n4727, n4728, n4729, n4731, n4732,
         n4733, n4734, n4735, n4737, n4740, n4743, n4744, n4745, n4746, n4747,
         n4749, n4750, n4751, n4752, n4753, n4755, n4758, n4761, n4762, n4763,
         n4764, n4765, n4767, n4768, n4769, n4770, n4771, n4773, n4776, n4779,
         n4780, n4781, n4782, n4783, n4785, n4786, n4787, n4788, n4789, n4791,
         n4794, n4797, n4798, n4799, n4800, n4801, n4803, n4804, n4805, n4806,
         n4807, n4809, n4812, n4815, n4816, n4817, n4818, n4819, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4840, n4843, n4844, n4847,
         n4848, n4849, n4853, n4854, n4857, n4858, n4859, n4860, n4861, n4866,
         n4867, n4870, n4871, n4872, n4873, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, N34665, N34664, N34663, N34662,
         N34661, N34660, N34659, N34658, N34657, N34656, N34655, N34654,
         N34653, N34652, N34651, N34650, N34649, N34648, N34647, N34646,
         N34645, N34644, N34643, N34642, N34641, N34640, N34639, N34638,
         N34637, N34636, N34635, N34634, N34633, N34632, N34631, N34630,
         N34629, N34628, N34627, N34626, N34625, N34624, N34623, N34622,
         N34621, N34620, N34619, N34618, N34617, N34616, N34615, N34614,
         N34613, N34612, N34611, N34610, N34609, N34608, N34607, N34606,
         N34605, N34604, N34603, N34602, N34601, N34600, N34599, N34598,
         N34597, N34596, N34595, N34594, N34593, N34592, N34591, N34590,
         N34589, N34588, N34587, N34586, N34585, N34584, N34583, N34582,
         N34581, N34580, N34579, N34578, N34577, N34576, N34575, N34574,
         N34573, N34572, N34571, N34570, N34569, N34568, N34567, N34566,
         N34565, N34564, N34563, N34562, N34561, N34560, N34559, N34558,
         N34557, N34556, N34555, N34554, N34553, N34552, N34551, N34550,
         N34549, N34548, N34547, N34546, N34545, N34544, N34543, N34542,
         N34541, N34540, N34539, N34537, N34536, N34535, N34534, N34533,
         N34532, N34531, N34530, N34529, N34528, N34527, N34526, N34525,
         N34524, N34523, N34522, N34521, N34520, N34519, N34518, N34517,
         N34516, N34515, N34514, N34513, N34512, N34511, N34510, N34509,
         N34508, N34507, N34506, N34505, N34504, N34503, N34502, N34501,
         N34500, N34499, N34498, N34497, N34496, N34495, N34494, N34493,
         N34492, N34491, N34490, N34489, N34488, N34487, N34486, N34485,
         N34484, N34483, N34482, N34481, N34480, N34479, N34478, N34477,
         N34476, N34475, N34474, N34473, N34472, N34471, N34470, N34469,
         N34468, N34467, N34466, N34465, N34464, N34463, N34462, N34461,
         N34460, N34459, N34458, N34457, N34456, N34455, N34454, N34453,
         N34452, N34451, N34450, N34449, N34448, N34447, N34446, N34445,
         N34444, N34443, N34442, N34441, N34440, N34439, N34438, N34437,
         N34436, N34435, N34434, N34433, N34432, N34431, N34430, N34429,
         N34428, N34427, N34426, N34425, N34424, N34423, N34422, N34421,
         N34420, N34419, N34418, N34417, N34416, N34415, N34414, N34413,
         N34412, N34411, N34410, N34409, N34408, N34407, N34406, N34405,
         N34404, N34403, N34402, N34401, N34400, N34399, N34398, N34397,
         N34396, N34395, N34394, N34393, N34392, N34391, N34390, N34389,
         N34388, N34387, N34386, N34385, N34384, N34383, N34382, N34381,
         N34380, N34379, N34378, N34377, N34376, N34375, N34374, N34373,
         N34372, N34371, N34370, N34369, N34368, N34367, N34366, N34365,
         N34364, N34363, N34362, N34361, N34360, N34359, N34358, N34357,
         N34356, N34355, N34354, N34353, N34352, N34351, N34350, N34349,
         N34348, N34347, N34345, N34344, N34343, N34342, N34341, N34340,
         N34339, N34338, N34337, N34336, N34335, N34334, N34333, N34332,
         N34331, N34330, N34329, N34328, N34327, N34326, N34325, N34324,
         N34323, N34322, N34321, N34320, N34319, N34318, N34317, N34316,
         N34315, N34314, N34313, N34312, N34311, N34310, N34309, N34308,
         N34307, N34306, N34305, N34304, N34303, N34302, N34301, N34300,
         N34299, N34298, N34297, N34296, N34295, N34294, N34293, N34292,
         N34291, N34290, N34289, N34288, N34287, N34286, N34285, N34284,
         N34283, N34282, N34281, N34280, N34279, N34278, N34277, N34276,
         N34275, N34274, N34273, N34272, N34271, N34270, N34269, N34268,
         N34267, N34266, N34265, N34264, N34263, N34262, N34261, N34260,
         N34259, N34258, N34257, N34256, N34255, N34254, N34253, N34252,
         N34251, N34250, N34249, N34248, N34247, N34246, N34245, N34244,
         N34243, N34242, N34241, N34240, N34239, N34238, N34237, N34236,
         N34235, N34234, N34233, N34232, N34231, N34230, N34229, N34228,
         N34227, N34226, N34225, N34224, N34223, N34222, N34221, N34220,
         N34219, N34217, N34216, N34215, N34214, N34213, N34212, N34211,
         N34210, N34209, N34208, N34207, N34206, N34205, N34204, N34203,
         N34202, N34201, N34200, N34199, N34198, N34197, N34196, N34195,
         N34194, N34193, N34192, N34191, N34190, N34189, N34188, N34187,
         N34186, N34185, N34184, N34183, N34182, N34181, N34180, N34179,
         N34178, N34177, N34176, N34175, N34174, N34173, N34172, N34171,
         N34170, N34169, N34168, N34167, N34166, N34165, N34164, N34163,
         N34162, N34161, N34160, N34159, N34158, N34157, N34156, N34155,
         N34153, N34152, N34151, N34150, N34149, N34148, N34147, N34146,
         N34145, N34144, N34143, N34142, N34141, N34140, N34139, N34138,
         N34137, N34136, N34135, N34134, N34133, N34132, N34131, N34130,
         N34129, N34128, N34127, N34126, N34125, N34124, N34123, N34122,
         N34121, N34120, N34119, N34118, N34117, N34116, N34115, N34114,
         N34113, N34112, N34111, N34110, N34109, N34108, N34107, N34106,
         N34105, N34104, N34103, N34102, N34101, N34100, N34099, N34098,
         N34097, N34096, N34095, N34094, N34093, N34092, N34091, N34090,
         N31273, N31272, N31271, N31270, N31269, N31268, N31267, N31266,
         N31265, N31264, N31263, N31262, N31261, N31260, N31259, N31258,
         N31257, N31256, N31255, N31254, N31253, N31252, N31251, N31250,
         N31249, N31248, N31247, N31246, N31245, N31244, N31243, N31242,
         N31241, N31240, N31239, N31238, N31237, N31236, N31235, N31234,
         N31233, N31232, N31231, N31230, N31229, N31228, N31227, N31226,
         N31225, N31224, N31223, N31222, N31221, N31220, N31219, N31218,
         N31217, N31216, N31215, N31214, N31213, N31212, N31211, N31210,
         N31209, N31208, N31207, N31206, N31205, N31204, N31203, N31202,
         N31201, N31200, N31199, N31198, N31197, N31196, N31195, N31194,
         N31193, N31192, N31191, N31190, N31189, N31188, N31187, N31186,
         N31185, N31184, N31183, N31182, N31181, N31180, N31179, N31178,
         N31177, N31176, N31175, N31174, N31173, N31172, N31171, N31170,
         N31169, N31168, N31167, N31166, N31165, N31164, N31163, N31162,
         N31161, N31160, N31159, N31158, N31157, N31156, N31155, N31154,
         N31153, N31152, N31151, N31150, N31149, N31148, N31147, N31145,
         N31144, N31143, N31142, N31141, N31140, N31139, N31138, N31137,
         N31136, N31135, N31134, N31133, N31132, N31131, N31130, N31129,
         N31128, N31127, N31126, N31125, N31124, N31123, N31122, N31121,
         N31120, N31119, N31118, N31117, N31116, N31115, N31114, N31113,
         N31112, N31111, N31110, N31109, N31108, N31107, N31106, N31105,
         N31104, N31103, N31102, N31101, N31100, N31099, N31098, N31097,
         N31096, N31095, N31094, N31093, N31092, N31091, N31090, N31089,
         N31088, N31087, N31086, N31085, N31084, N31083, N31082, N31081,
         N31080, N31079, N31078, N31077, N31076, N31075, N31074, N31073,
         N31072, N31071, N31070, N31069, N31068, N31067, N31066, N31065,
         N31064, N31063, N31062, N31061, N31060, N31059, N31058, N31057,
         N31056, N31055, N31054, N31053, N31052, N31051, N31050, N31049,
         N31048, N31047, N31046, N31045, N31044, N31043, N31042, N31041,
         N31040, N31039, N31038, N31037, N31036, N31035, N31034, N31033,
         N31032, N31031, N31030, N31029, N31028, N31027, N31026, N31025,
         N31024, N31023, N31022, N31021, N31020, N31019, N31018, N31017,
         N31016, N31015, N31014, N31013, N31012, N31011, N31010, N31009,
         N31008, N31007, N31006, N31005, N31004, N31003, N31002, N31001,
         N31000, N30999, N30998, N30997, N30996, N30995, N30994, N30993,
         N30992, N30991, N30990, N30989, N30988, N30987, N30986, N30985,
         N30984, N30983, N30982, N30981, N30980, N30979, N30978, N30977,
         N30976, N30975, N30974, N30973, N30972, N30971, N30970, N30969,
         N30968, N30967, N30966, N30965, N30964, N30963, N30962, N30961,
         N30960, N30959, N30958, N30957, N30956, N30955, N30953, N30952,
         N30951, N30950, N30949, N30948, N30947, N30946, N30945, N30944,
         N30943, N30942, N30941, N30940, N30939, N30938, N30937, N30936,
         N30935, N30934, N30933, N30932, N30931, N30930, N30929, N30928,
         N30927, N30926, N30925, N30924, N30923, N30922, N30921, N30920,
         N30919, N30918, N30917, N30916, N30915, N30914, N30913, N30912,
         N30911, N30910, N30909, N30908, N30907, N30906, N30905, N30904,
         N30903, N30902, N30901, N30900, N30899, N30898, N30897, N30896,
         N30895, N30894, N30893, N30892, N30891, N30890, N30889, N30888,
         N30887, N30886, N30885, N30884, N30883, N30882, N30881, N30880,
         N30879, N30878, N30877, N30876, N30875, N30874, N30873, N30872,
         N30871, N30870, N30869, N30868, N30867, N30866, N30865, N30864,
         N30863, N30862, N30861, N30860, N30859, N30858, N30857, N30856,
         N30855, N30854, N30853, N30852, N30851, N30850, N30849, N30848,
         N30847, N30846, N30845, N30844, N30843, N30842, N30841, N30840,
         N30839, N30838, N30837, N30836, N30835, N30834, N30833, N30832,
         N30831, N30830, N30829, N30828, N30827, N30826, N30825, N30824,
         N30823, N30822, N30821, N30820, N30819, N30818, N30817, N30816,
         N30815, N30814, N30813, N30812, N30811, N30810, N30809, N30808,
         N30807, N30806, N30805, N30804, N30803, N30802, N30801, N30800,
         N30799, N30798, N30797, N30796, N30795, N30794, N30793, N30792,
         N30791, N30790, N30789, N30788, N30787, N30786, N30785, N30784,
         N30783, N30782, N30781, N30780, N30779, N30778, N30777, N30776,
         N30775, N30774, N30773, N30772, N30771, N30770, N30769, N30768,
         N30767, N30766, N30765, N30764, N30763, N30313, N30312, N30311,
         N30310, N30309, N30308, N30307, N30306, N30305, N30304, N30303,
         N30302, N30301, N30300, N30299, N30298, N30297, N30296, N30295,
         N30294, N30293, N30292, N30291, N30290, N30289, N30288, N30287,
         N30286, N30285, N30284, N30283, N30282, N30281, N30280, N30279,
         N30278, N30277, N30276, N30275, N30274, N30273, N30272, N30271,
         N30270, N30269, N30268, N30267, N30266, N30265, N30264, N30263,
         N30262, N30261, N30260, N30259, N30258, N30257, N30256, N30255,
         N30254, N30253, N30252, N30251, N30250, N30249, N30248, N30247,
         N30246, N30245, N30244, N30243, N30242, N30241, N30240, N30239,
         N30238, N30237, N30236, N30235, N30234, N30233, N30232, N30231,
         N30230, N30229, N30228, N30227, N30226, N30225, N30224, N30223,
         N30222, N30221, N30220, N30219, N30218, N30217, N30216, N30215,
         N30214, N30213, N30212, N30211, N30210, N30209, N30208, N30207,
         N30206, N30205, N30204, N30203, N30202, N30201, N30200, N30199,
         N30198, N30197, N30196, N30195, N30194, N30193, N30192, N30191,
         N30190, N30189, N30188, N30187, N30185, N30184, N30183, N30182,
         N30181, N30180, N30179, N30178, N30177, N30176, N30175, N30174,
         N30173, N30172, N30171, N30170, N30169, N30168, N30167, N30166,
         N30165, N30164, N30163, N30162, N30161, N30160, N30159, N30158,
         N30157, N30156, N30155, N30154, N30153, N30152, N30151, N30150,
         N30149, N30148, N30147, N30146, N30145, N30144, N30143, N30142,
         N30141, N30140, N30139, N30138, N30137, N30136, N30135, N30134,
         N30133, N30132, N30131, N30130, N30129, N30128, N30127, N30126,
         N30125, N30124, N30123, N30122, N30121, N30120, N30119, N30118,
         N30117, N30116, N30115, N30114, N30113, N30112, N30111, N30110,
         N30109, N30108, N30107, N30106, N30105, N30104, N30103, N30102,
         N30101, N30100, N30099, N30098, N30097, N30096, N30095, N30094,
         N30093, N30092, N30091, N30090, N30089, N30088, N30087, N30086,
         N30085, N30084, N30083, N30082, N30081, N30080, N30079, N30078,
         N30077, N30076, N30075, N30074, N30073, N30072, N30071, N30070,
         N30069, N30068, N30067, N30066, N30065, N30064, N30063, N30062,
         N30061, N30060, N30059, N30058, N30057, N30056, N30055, N30054,
         N30053, N30052, N30051, N30050, N30049, N30048, N30047, N30046,
         N30045, N30044, N30043, N30042, N30041, N30040, N30039, N30038,
         N30037, N30036, N30035, N30034, N30033, N30032, N30031, N30030,
         N30029, N30028, N30027, N30026, N30025, N30024, N30023, N30022,
         N30021, N30020, N30019, N30018, N30017, N30016, N30015, N30014,
         N30013, N30012, N30011, N30010, N30009, N30008, N30007, N30006,
         N30005, N30004, N30003, N30002, N30001, N30000, N29999, N29998,
         N29997, N29996, N29995, N29993, N29992, N29991, N29990, N29989,
         N29988, N29987, N29986, N29985, N29984, N29983, N29982, N29981,
         N29980, N29979, N29978, N29977, N29976, N29975, N29974, N29973,
         N29972, N29971, N29970, N29969, N29968, N29967, N29966, N29965,
         N29964, N29963, N29962, N29961, N29960, N29959, N29958, N29957,
         N29956, N29955, N29954, N29953, N29952, N29951, N29950, N29949,
         N29948, N29947, N29946, N29945, N29944, N29943, N29942, N29941,
         N29940, N29939, N29938, N29937, N29936, N29935, N29934, N29933,
         N29932, N29931, N29930, N33577, N33576, N33575, N33574, N33573,
         N33572, N33571, N33570, N33569, N33568, N33567, N33566, N33565,
         N33564, N33563, N33562, N33561, N33560, N33559, N33558, N33557,
         N33556, N33555, N33554, N33553, N33552, N33551, N33550, N33549,
         N33548, N33547, N33546, N33545, N33544, N33543, N33542, N33541,
         N33540, N33539, N33538, N33537, N33536, N33535, N33534, N33533,
         N33532, N33531, N33530, N33529, N33528, N33527, N33526, N33525,
         N33524, N33523, N33522, N33521, N33520, N33519, N33518, N33517,
         N33516, N33515, N33513, N33512, N33511, N33510, N33509, N33508,
         N33507, N33506, N33505, N33504, N33503, N33502, N33501, N33500,
         N33499, N33498, N33497, N33496, N33495, N33494, N33493, N33492,
         N33491, N33490, N33489, N33488, N33487, N33486, N33485, N33484,
         N33483, N33482, N33481, N33480, N33479, N33478, N33477, N33476,
         N33475, N33474, N33473, N33472, N33471, N33470, N33469, N33468,
         N33467, N33466, N33465, N33464, N33463, N33462, N33461, N33460,
         N33459, N33458, N33457, N33456, N33455, N33454, N33453, N33452,
         N33451, N33450, N33449, N33448, N33447, N33446, N33445, N33444,
         N33443, N33442, N33441, N33440, N33439, N33438, N33437, N33436,
         N33435, N33434, N33433, N33432, N33431, N33430, N33429, N33428,
         N33427, N33426, N33425, N33424, N33423, N33422, N33421, N33420,
         N33419, N33418, N33417, N33416, N33415, N33414, N33413, N33412,
         N33411, N33410, N33409, N33408, N33407, N33406, N33405, N33404,
         N33403, N33402, N33401, N33400, N33399, N33398, N33397, N33396,
         N33395, N33394, N33393, N33392, N33391, N33390, N33389, N33388,
         N33387, N33386, N33385, N33384, N33383, N33382, N33381, N33380,
         N33379, N33378, N33377, N33376, N33375, N33374, N33373, N33372,
         N33371, N33370, N33369, N33368, N33367, N33366, N33365, N33364,
         N33363, N33362, N33361, N33360, N33359, N33358, N33357, N33356,
         N33355, N33354, N33353, N33352, N33351, N33350, N33349, N33348,
         N33347, N33346, N33345, N33344, N33343, N33342, N33341, N33340,
         N33339, N33338, N33337, N33336, N33335, N33334, N33333, N33332,
         N33331, N33330, N33329, N33328, N33327, N33326, N33325, N33324,
         N33323, N33322, N33321, N33320, N33319, N33318, N33317, N33316,
         N33315, N33314, N33313, N33312, N33311, N33310, N33309, N33308,
         N33307, N33306, N33305, N33304, N33303, N33302, N33301, N33300,
         N33299, N33298, N33297, N33296, N33295, N33294, N33293, N33292,
         N33291, N33290, N33289, N33288, N33287, N33286, N33285, N33284,
         N33283, N33282, N33281, N33280, N33279, N33278, N33277, N33276,
         N33275, N33274, N33273, N33272, N33271, N33270, N33269, N33268,
         N33267, N33266, N33265, N33264, N33263, N33262, N33261, N33260,
         N33259, N33258, N33257, N33256, N33255, N33254, N33253, N33252,
         N33251, N33250, N33249, N33248, N33247, N33246, N33245, N33244,
         N33243, N33242, N33241, N33240, N33239, N33238, N33237, N33236,
         N33235, N33234, N33233, N33232, N33231, N33230, N33229, N33228,
         N33227, N33226, N33225, N33224, N33223, N33222, N33221, N33220,
         N33219, N33218, N33217, N33216, N33215, N33214, N33213, N33212,
         N33211, N33210, N33209, N33208, N33207, N33206, N33205, N33204,
         N33203, N33202, N33201, N33200, N33199, N33198, N33197, N33196,
         N33195, N33193, N33192, N33191, N33190, N33189, N33188, N33187,
         N33186, N33185, N33184, N33183, N33182, N33181, N33180, N33179,
         N33178, N33177, N33176, N33175, N33174, N33173, N33172, N33171,
         N33170, N33169, N33168, N33167, N33166, N33165, N33164, N33163,
         N33162, N33161, N33160, N33159, N33158, N33157, N33156, N33155,
         N33154, N33153, N33152, N33151, N33150, N33149, N33148, N33147,
         N33146, N33145, N33144, N33143, N33142, N33141, N33140, N33139,
         N33138, N33137, N33136, N33135, N33134, N33133, N33132, N33131,
         N33129, N33128, N33127, N33126, N33125, N33124, N33123, N33122,
         N33121, N33120, N33119, N33118, N33117, N33116, N33115, N33114,
         N33113, N33112, N33111, N33110, N33109, N33108, N33107, N33106,
         N33105, N33104, N33103, N33102, N33101, N33100, N33099, N33098,
         N33097, N33096, N33095, N33094, N33093, N33092, N33091, N33090,
         N33089, N33088, N33087, N33086, N33085, N33084, N33083, N33082,
         N33081, N33080, N33079, N33078, N33077, N33076, N33075, N33074,
         N33073, N33072, N33071, N33070, N33069, N33068, N33067, N32617,
         N32616, N32615, N32614, N32613, N32612, N32611, N32610, N32609,
         N32608, N32607, N32606, N32605, N32604, N32603, N32602, N32601,
         N32600, N32599, N32598, N32597, N32596, N32595, N32594, N32593,
         N32592, N32591, N32590, N32589, N32588, N32587, N32586, N32585,
         N32584, N32583, N32582, N32581, N32580, N32579, N32578, N32577,
         N32576, N32575, N32574, N32573, N32572, N32571, N32570, N32569,
         N32568, N32567, N32566, N32565, N32564, N32563, N32562, N32561,
         N32560, N32559, N32558, N32557, N32556, N32555, N32554, N32553,
         N32552, N32551, N32550, N32549, N32548, N32547, N32546, N32545,
         N32544, N32543, N32542, N32541, N32540, N32539, N32538, N32537,
         N32536, N32535, N32534, N32533, N32532, N32531, N32530, N32529,
         N32528, N32527, N32526, N32525, N32524, N32523, N32522, N32521,
         N32520, N32519, N32518, N32517, N32516, N32515, N32514, N32513,
         N32512, N32511, N32510, N32509, N32508, N32507, N32506, N32505,
         N32504, N32503, N32502, N32501, N32500, N32499, N32498, N32497,
         N32496, N32495, N32494, N32493, N32492, N32491, N32490, N32489,
         N32488, N32487, N32486, N32485, N32484, N32483, N32482, N32481,
         N32480, N32479, N32478, N32477, N32476, N32475, N32474, N32473,
         N32472, N32471, N32470, N32469, N32468, N32467, N32466, N32465,
         N32464, N32463, N32462, N32461, N32460, N32459, N32458, N32457,
         N32456, N32455, N32454, N32453, N32452, N32451, N32450, N32449,
         N32448, N32447, N32446, N32445, N32444, N32443, N32442, N32441,
         N32440, N32439, N32438, N32437, N32436, N32435, N32434, N32433,
         N32432, N32431, N32430, N32429, N32428, N32427, N32426, N32425,
         N32424, N32423, N32422, N32421, N32420, N32419, N32418, N32417,
         N32416, N32415, N32414, N32413, N32412, N32411, N32410, N32409,
         N32408, N32407, N32406, N32405, N32404, N32403, N32402, N32401,
         N32400, N32399, N32398, N32397, N32396, N32395, N32394, N32393,
         N32392, N32391, N32390, N32389, N32388, N32387, N32386, N32385,
         N32384, N32383, N32382, N32381, N32380, N32379, N32378, N32377,
         N32376, N32375, N32374, N32373, N32372, N32371, N32370, N32369,
         N32368, N32367, N32366, N32365, N32364, N32363, N32362, N32361,
         N32360, N32359, N32358, N32357, N32356, N32355, N32354, N32353,
         N32352, N32351, N32350, N32349, N32348, N32347, N32346, N32345,
         N32344, N32343, N32342, N32341, N32340, N32339, N32338, N32337,
         N32336, N32335, N32334, N32333, N32332, N32331, N32330, N32329,
         N32328, N32327, N32326, N32325, N32324, N32323, N32322, N32321,
         N32320, N32319, N32318, N32317, N32316, N32315, N32314, N32313,
         N32312, N32311, N32310, N32309, N32308, N32307, N32306, N32305,
         N32304, N32303, N32302, N32301, N32300, N32299, N32297, N32296,
         N32295, N32294, N32293, N32292, N32291, N32290, N32289, N32288,
         N32287, N32286, N32285, N32284, N32283, N32282, N32281, N32280,
         N32279, N32278, N32277, N32276, N32275, N32274, N32273, N32272,
         N32271, N32270, N32269, N32268, N32267, N32266, N32265, N32264,
         N32263, N32262, N32261, N32260, N32259, N32258, N32257, N32256,
         N32255, N32254, N32253, N32252, N32251, N32250, N32249, N32248,
         N32247, N32246, N32245, N32244, N32243, N32242, N32241, N32240,
         N32239, N32238, N32237, N32236, N32235, N31849, N31848, N31847,
         N31846, N31845, N31844, N31843, N31842, N31841, N31840, N31839,
         N31838, N31837, N31836, N31835, N31834, N31833, N31832, N31831,
         N31830, N31829, N31828, N31827, N31826, N31825, N31824, N31823,
         N31822, N31821, N31820, N31819, N31818, N31817, N31816, N31815,
         N31814, N31813, N31812, N31811, N31810, N31809, N31808, N31807,
         N31806, N31805, N31804, N31803, N31802, N31801, N31800, N31799,
         N31798, N31797, N31796, N31795, N31794, N31793, N31792, N31791,
         N31790, N31789, N31788, N31787, N31786, N31785, N31784, N31783,
         N31782, N31781, N31780, N31779, N31778, N31777, N31776, N31775,
         N31774, N31773, N31772, N31771, N31770, N31769, N31768, N31767,
         N31766, N31765, N31764, N31763, N31762, N31761, N31760, N31759,
         N31758, N31757, N31756, N31755, N31754, N31753, N31752, N31751,
         N31750, N31749, N31748, N31747, N31746, N31745, N31744, N31743,
         N31742, N31741, N31740, N31739, N31738, N31737, N31736, N31735,
         N31734, N31733, N31732, N31731, N31730, N31729, N31728, N31727,
         N31726, N31725, N31724, N31723, N31721, N31720, N31719, N31718,
         N31717, N31716, N31715, N31714, N31713, N31712, N31711, N31710,
         N31709, N31708, N31707, N31706, N31705, N31704, N31703, N31702,
         N31701, N31700, N31699, N31698, N31697, N31696, N31695, N31694,
         N31693, N31692, N31691, N31690, N31689, N31688, N31687, N31686,
         N31685, N31684, N31683, N31682, N31681, N31680, N31679, N31678,
         N31677, N31676, N31675, N31674, N31673, N31672, N31671, N31670,
         N31669, N31668, N31667, N31666, N31665, N31664, N31663, N31662,
         N31661, N31660, N31659, N31657, N31656, N31655, N31654, N31653,
         N31652, N31651, N31650, N31649, N31648, N31647, N31646, N31645,
         N31644, N31643, N31642, N31641, N31640, N31639, N31638, N31637,
         N31636, N31635, N31634, N31633, N31632, N31631, N31630, N31629,
         N31628, N31627, N31626, N31625, N31624, N31623, N31622, N31621,
         N31620, N31619, N31618, N31617, N31616, N31615, N31614, N31613,
         N31612, N31611, N31610, N31609, N31608, N31607, N31606, N31605,
         N31604, N31603, N31602, N31601, N31600, N31599, N31598, N31597,
         N31596, N31595, N31594, N29545, N29544, N29543, N29542, N29541,
         N29540, N29539, N29538, N29537, N29536, N29535, N29534, N29533,
         N29532, N29531, N29530, N29529, N29528, N29527, N29526, N29525,
         N29524, N29523, N29522, N29521, N29520, N29519, N29518, N29517,
         N29516, N29515, N29514, N29513, N29512, N29511, N29510, N29509,
         N29508, N29507, N29506, N29505, N29504, N29503, N29502, N29501,
         N29500, N29499, N29498, N29497, N29496, N29495, N29494, N29493,
         N29492, N29491, N29490, N29489, N29488, N29487, N29486, N29485,
         N29484, N29483, N29481, N29480, N29479, N29478, N29477, N29476,
         N29475, N29474, N29473, N29472, N29471, N29470, N29469, N29468,
         N29467, N29466, N29465, N29464, N29463, N29462, N29461, N29460,
         N29459, N29458, N29457, N29456, N29455, N29454, N29453, N29452,
         N29451, N29450, N29449, N29448, N29447, N29446, N29445, N29444,
         N29443, N29442, N29441, N29440, N29439, N29438, N29437, N29436,
         N29435, N29434, N29433, N29432, N29431, N29430, N29429, N29428,
         N29427, N29426, N29425, N29424, N29423, N29422, N29421, N29420,
         N29419, N29417, N29416, N29415, N29414, N29413, N29412, N29411,
         N29410, N29409, N29408, N29407, N29406, N29405, N29404, N29403,
         N29402, N29401, N29400, N29399, N29398, N29397, N29396, N29395,
         N29394, N29393, N29392, N29391, N29390, N29389, N29388, N29387,
         N29386, N29385, N29384, N29383, N29382, N29381, N29380, N29379,
         N29378, N29377, N29376, N29375, N29374, N29373, N29372, N29371,
         N29370, N29369, N29368, N29367, N29366, N29365, N29364, N29363,
         N29362, N29361, N29360, N29359, N29358, N29357, N29356, N29355,
         N29354, N29353, N29352, N29351, N29350, N29349, N29348, N29347,
         N29346, N29345, N29344, N29343, N29342, N29341, N29340, N29339,
         N29338, N29337, N29336, N29335, N29334, N29333, N29332, N29331,
         N29330, N29329, N29328, N29327, N29326, N29325, N29324, N29323,
         N29322, N29321, N29320, N29319, N29318, N29317, N29316, N29315,
         N29314, N29313, N29312, N29311, N29310, N29309, N29308, N29307,
         N29306, N29305, N29304, N29303, N29302, N29301, N29300, N29299,
         N29298, N29297, N29296, N29295, N29294, N29293, N29292, N29291,
         N29290, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6627, n6629, n6631, n6633, n6635, n6637,
         n6639, n6641, n6643, n6645, n6647, n6649, n6651, n6653, n6655, n6657,
         n6659, n6661, n6663, n6665, n6667, n6669, n6671, n6673, n6675, n6677,
         n6679, n6681, n6683, n6685, n6687, n6689, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398;
  wire   [31:0] inCount;
  wire   [1:0] state;
  wire   [31:0] xCount;
  wire   [31:0] iCount;
  wire   [1:0] state_next;
  wire   [31:0] outCount_next;
  wire   [31:0] outCount;
  wire   [31:0] xCount_next;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120;
  assign N2348 = b_in[15];
  assign N35189 = in_en;

  OAI221X2 U1380 ( .A0(n8315), .A1(n279), .B0(n7719), .B1(n277), .C0(n787), 
        .Y(N34024) );
  OAI221X2 U1384 ( .A0(n8315), .A1(n287), .B0(n7719), .B1(n285), .C0(n790), 
        .Y(N34023) );
  OAI221X2 U1388 ( .A0(n8315), .A1(n295), .B0(n7719), .B1(n293), .C0(n793), 
        .Y(N34022) );
  OAI221X2 U1392 ( .A0(n8315), .A1(n303), .B0(n7719), .B1(n301), .C0(n796), 
        .Y(N34021) );
  OAI221X2 U1396 ( .A0(n8315), .A1(n311), .B0(n7719), .B1(n309), .C0(n799), 
        .Y(N34020) );
  OAI221X2 U1400 ( .A0(n8315), .A1(n319), .B0(n7719), .B1(n317), .C0(n802), 
        .Y(N34019) );
  OAI221X2 U1404 ( .A0(n8315), .A1(n327), .B0(n7719), .B1(n325), .C0(n805), 
        .Y(N34018) );
  OAI221X2 U1408 ( .A0(n8315), .A1(n335), .B0(n7719), .B1(n333), .C0(n808), 
        .Y(N34017) );
  OAI221X2 U1412 ( .A0(n8315), .A1(n343), .B0(n7719), .B1(n341), .C0(n811), 
        .Y(N34016) );
  OAI221X2 U1416 ( .A0(n8315), .A1(n351), .B0(n7719), .B1(n349), .C0(n814), 
        .Y(N34015) );
  OAI221X2 U1420 ( .A0(n8315), .A1(n359), .B0(n7719), .B1(n357), .C0(n817), 
        .Y(N34014) );
  OAI221X2 U1424 ( .A0(n8323), .A1(n367), .B0(n7720), .B1(n365), .C0(n820), 
        .Y(N34013) );
  OAI221X2 U1428 ( .A0(n8323), .A1(n375), .B0(n7720), .B1(n373), .C0(n823), 
        .Y(N34012) );
  OAI221X2 U1432 ( .A0(n8323), .A1(n383), .B0(n7720), .B1(n381), .C0(n826), 
        .Y(N34011) );
  OAI221X2 U1436 ( .A0(n8323), .A1(n391), .B0(n7720), .B1(n389), .C0(n829), 
        .Y(N34010) );
  OAI221X2 U1440 ( .A0(n8323), .A1(n399), .B0(n7720), .B1(n397), .C0(n832), 
        .Y(N34009) );
  OAI221X2 U1444 ( .A0(n8323), .A1(n407), .B0(n7720), .B1(n405), .C0(n835), 
        .Y(N34008) );
  OAI221X2 U1448 ( .A0(n8323), .A1(n415), .B0(n7720), .B1(n413), .C0(n838), 
        .Y(N34007) );
  OAI221X2 U1452 ( .A0(n8323), .A1(n423), .B0(n7720), .B1(n421), .C0(n841), 
        .Y(N34006) );
  OAI221X2 U1456 ( .A0(n8323), .A1(n431), .B0(n7720), .B1(n429), .C0(n844), 
        .Y(N34005) );
  OAI221X2 U1460 ( .A0(n8323), .A1(n439), .B0(n7720), .B1(n437), .C0(n847), 
        .Y(N34004) );
  OAI221X2 U1464 ( .A0(n8319), .A1(n447), .B0(n7720), .B1(n445), .C0(n850), 
        .Y(N34003) );
  OAI221X2 U1468 ( .A0(n8319), .A1(n455), .B0(n7720), .B1(n453), .C0(n853), 
        .Y(N34002) );
  OAI221X2 U1472 ( .A0(n8319), .A1(n463), .B0(n7720), .B1(n461), .C0(n856), 
        .Y(N34001) );
  OAI221X2 U1476 ( .A0(n8314), .A1(n471), .B0(n7721), .B1(n469), .C0(n859), 
        .Y(N34000) );
  OAI221X2 U1480 ( .A0(n8314), .A1(n479), .B0(n7721), .B1(n477), .C0(n862), 
        .Y(N33999) );
  OAI221X2 U1484 ( .A0(n8309), .A1(n487), .B0(n7721), .B1(n485), .C0(n865), 
        .Y(N33998) );
  OAI221X2 U1488 ( .A0(n8314), .A1(n495), .B0(n7721), .B1(n493), .C0(n868), 
        .Y(N33997) );
  OAI221X2 U1492 ( .A0(n8314), .A1(n503), .B0(n7721), .B1(n501), .C0(n871), 
        .Y(N33996) );
  OAI221X2 U1496 ( .A0(n8307), .A1(n511), .B0(n7721), .B1(n509), .C0(n874), 
        .Y(N33995) );
  OAI221X2 U1500 ( .A0(n8317), .A1(n519), .B0(n7721), .B1(n517), .C0(n877), 
        .Y(N33994) );
  OAI221X2 U1504 ( .A0(n8318), .A1(n527), .B0(n7721), .B1(n525), .C0(n880), 
        .Y(N33993) );
  OAI221X2 U1508 ( .A0(n8314), .A1(n535), .B0(n7721), .B1(n533), .C0(n883), 
        .Y(N33992) );
  OAI221X2 U1512 ( .A0(n8309), .A1(n543), .B0(n7721), .B1(n541), .C0(n886), 
        .Y(N33991) );
  OAI221X2 U1516 ( .A0(n8314), .A1(n551), .B0(n7721), .B1(n549), .C0(n889), 
        .Y(N33990) );
  OAI221X2 U1520 ( .A0(n8312), .A1(n559), .B0(n7721), .B1(n557), .C0(n892), 
        .Y(N33989) );
  OAI221X2 U1524 ( .A0(n8315), .A1(n567), .B0(n7721), .B1(n565), .C0(n895), 
        .Y(N33988) );
  OAI221X2 U1528 ( .A0(n8315), .A1(n575), .B0(n7722), .B1(n573), .C0(n898), 
        .Y(N33987) );
  OAI221X2 U1532 ( .A0(n8316), .A1(n583), .B0(n7722), .B1(n581), .C0(n901), 
        .Y(N33986) );
  OAI221X2 U1536 ( .A0(n8316), .A1(n591), .B0(n7722), .B1(n589), .C0(n904), 
        .Y(N33985) );
  OAI221X2 U1540 ( .A0(n8316), .A1(n599), .B0(n7722), .B1(n597), .C0(n907), 
        .Y(N33984) );
  OAI221X2 U1544 ( .A0(n8316), .A1(n607), .B0(n7722), .B1(n605), .C0(n910), 
        .Y(N33983) );
  OAI221X2 U1548 ( .A0(n8316), .A1(n615), .B0(n7722), .B1(n613), .C0(n913), 
        .Y(N33982) );
  OAI221X2 U1552 ( .A0(n8316), .A1(n623), .B0(n7722), .B1(n621), .C0(n916), 
        .Y(N33981) );
  OAI221X2 U1556 ( .A0(n8316), .A1(n631), .B0(n7722), .B1(n629), .C0(n919), 
        .Y(N33980) );
  OAI221X2 U1560 ( .A0(n8316), .A1(n639), .B0(n7722), .B1(n637), .C0(n922), 
        .Y(N33979) );
  OAI221X2 U1564 ( .A0(n8316), .A1(n647), .B0(n7722), .B1(n645), .C0(n925), 
        .Y(N33978) );
  OAI221X2 U1568 ( .A0(n8316), .A1(n655), .B0(n7722), .B1(n653), .C0(n928), 
        .Y(N33977) );
  OAI221X2 U1572 ( .A0(n8316), .A1(n663), .B0(n7722), .B1(n661), .C0(n931), 
        .Y(N33976) );
  OAI221X2 U1576 ( .A0(n8316), .A1(n671), .B0(n7722), .B1(n669), .C0(n934), 
        .Y(N33975) );
  OAI221X2 U1580 ( .A0(n8316), .A1(n679), .B0(n7723), .B1(n677), .C0(n937), 
        .Y(N33974) );
  OAI221X2 U1584 ( .A0(n8317), .A1(n687), .B0(n7723), .B1(n685), .C0(n940), 
        .Y(N33973) );
  OAI221X2 U1588 ( .A0(n8317), .A1(n695), .B0(n7723), .B1(n693), .C0(n943), 
        .Y(N33972) );
  OAI221X2 U1592 ( .A0(n8317), .A1(n703), .B0(n7723), .B1(n701), .C0(n946), 
        .Y(N33971) );
  OAI221X2 U1596 ( .A0(n8317), .A1(n711), .B0(n7723), .B1(n709), .C0(n949), 
        .Y(N33970) );
  OAI221X2 U1600 ( .A0(n8317), .A1(n719), .B0(n7723), .B1(n717), .C0(n952), 
        .Y(N33969) );
  OAI221X2 U1604 ( .A0(n8317), .A1(n727), .B0(n7723), .B1(n725), .C0(n955), 
        .Y(N33968) );
  OAI221X2 U1608 ( .A0(n8317), .A1(n735), .B0(n7723), .B1(n733), .C0(n958), 
        .Y(N33967) );
  OAI221X2 U1612 ( .A0(n8317), .A1(n743), .B0(n7723), .B1(n741), .C0(n961), 
        .Y(N33966) );
  OAI221X2 U1632 ( .A0(n8317), .A1(n267), .B0(n7724), .B1(n784), .C0(n976), 
        .Y(N33961) );
  OAI221X2 U1638 ( .A0(n8320), .A1(n277), .B0(n7724), .B1(n788), .C0(n981), 
        .Y(N33960) );
  OAI221X2 U2016 ( .A0(n8312), .A1(n977), .B0(n7727), .B1(n1296), .C0(n1297), 
        .Y(N33897) );
  OAI221X2 U2020 ( .A0(n8309), .A1(n982), .B0(n7716), .B1(n1300), .C0(n1301), 
        .Y(N33896) );
  OAI221X2 U2276 ( .A0(n8312), .A1(n1300), .B0(n7716), .B1(n1302), .C0(n1555), 
        .Y(N33832) );
  OAI221X2 U2280 ( .A0(n8312), .A1(n1304), .B0(n7716), .B1(n1306), .C0(n1558), 
        .Y(N33831) );
  OAI221X2 U2284 ( .A0(n8312), .A1(n1308), .B0(n7716), .B1(n1310), .C0(n1561), 
        .Y(N33830) );
  OAI221X2 U2288 ( .A0(n8312), .A1(n1312), .B0(n7716), .B1(n1314), .C0(n1564), 
        .Y(N33829) );
  OAI221X2 U2292 ( .A0(n8312), .A1(n1316), .B0(n7716), .B1(n1318), .C0(n1567), 
        .Y(N33828) );
  OAI221X2 U2296 ( .A0(n8312), .A1(n1320), .B0(n7716), .B1(n1322), .C0(n1570), 
        .Y(N33827) );
  OAI221X2 U2300 ( .A0(n8312), .A1(n1324), .B0(n7716), .B1(n1326), .C0(n1573), 
        .Y(N33826) );
  OAI221X2 U2304 ( .A0(n8312), .A1(n1328), .B0(n7716), .B1(n1330), .C0(n1576), 
        .Y(N33825) );
  OAI221X2 U2308 ( .A0(n8312), .A1(n1332), .B0(n7716), .B1(n1334), .C0(n1579), 
        .Y(N33824) );
  OAI221X2 U2312 ( .A0(n8318), .A1(n1336), .B0(n7733), .B1(n1338), .C0(n1582), 
        .Y(N33823) );
  OAI221X2 U2316 ( .A0(n8311), .A1(n1340), .B0(n7733), .B1(n1342), .C0(n1585), 
        .Y(N33822) );
  OAI221X2 U2320 ( .A0(n8318), .A1(n1344), .B0(n7733), .B1(n1346), .C0(n1588), 
        .Y(N33821) );
  OAI221X2 U2324 ( .A0(n8311), .A1(n1348), .B0(n7733), .B1(n1350), .C0(n1591), 
        .Y(N33820) );
  OAI221X2 U2328 ( .A0(n8318), .A1(n1352), .B0(n7740), .B1(n1354), .C0(n1594), 
        .Y(N33819) );
  OAI221X2 U2332 ( .A0(n8311), .A1(n1356), .B0(n7711), .B1(n1358), .C0(n1597), 
        .Y(N33818) );
  OAI221X2 U2336 ( .A0(n8318), .A1(n1360), .B0(n7711), .B1(n1362), .C0(n1600), 
        .Y(N33817) );
  OAI221X2 U2340 ( .A0(n8318), .A1(n1364), .B0(n7726), .B1(n1366), .C0(n1603), 
        .Y(N33816) );
  OAI221X2 U2344 ( .A0(n8318), .A1(n1368), .B0(n7717), .B1(n1370), .C0(n1606), 
        .Y(N33815) );
  OAI221X2 U2348 ( .A0(n8308), .A1(n1372), .B0(n7722), .B1(n1374), .C0(n1609), 
        .Y(N33814) );
  OAI221X2 U2352 ( .A0(n8308), .A1(n1376), .B0(n7722), .B1(n1378), .C0(n1612), 
        .Y(N33813) );
  OAI221X2 U2356 ( .A0(n8308), .A1(n1380), .B0(n7737), .B1(n1382), .C0(n1615), 
        .Y(N33812) );
  OAI221X2 U2360 ( .A0(n8308), .A1(n1384), .B0(n7737), .B1(n1386), .C0(n1618), 
        .Y(N33811) );
  OAI221X2 U2364 ( .A0(n8312), .A1(n1388), .B0(n7711), .B1(n1390), .C0(n1621), 
        .Y(N33810) );
  OAI221X2 U2368 ( .A0(n8317), .A1(n1392), .B0(n7711), .B1(n1394), .C0(n1624), 
        .Y(N33809) );
  OAI221X2 U2372 ( .A0(n8312), .A1(n1396), .B0(n7740), .B1(n1398), .C0(n1627), 
        .Y(N33808) );
  OAI221X2 U2376 ( .A0(n8312), .A1(n1400), .B0(n7740), .B1(n1402), .C0(n1630), 
        .Y(N33807) );
  OAI221X2 U2380 ( .A0(n8315), .A1(n1404), .B0(n7740), .B1(n1406), .C0(n1633), 
        .Y(N33806) );
  OAI221X2 U2384 ( .A0(n8312), .A1(n1408), .B0(n7728), .B1(n1410), .C0(n1636), 
        .Y(N33805) );
  OAI221X2 U2388 ( .A0(n8312), .A1(n1412), .B0(n7728), .B1(n1414), .C0(n1639), 
        .Y(N33804) );
  OAI221X2 U2392 ( .A0(n8312), .A1(n1416), .B0(n7728), .B1(n1418), .C0(n1642), 
        .Y(N33803) );
  OAI221X2 U2396 ( .A0(n8311), .A1(n1420), .B0(n7728), .B1(n1422), .C0(n1645), 
        .Y(N33802) );
  OAI221X2 U2400 ( .A0(n8311), .A1(n1424), .B0(n7728), .B1(n1426), .C0(n1648), 
        .Y(N33801) );
  OAI221X2 U2404 ( .A0(n8318), .A1(n1428), .B0(n7726), .B1(n1430), .C0(n1651), 
        .Y(N33800) );
  OAI221X2 U2408 ( .A0(n8318), .A1(n1432), .B0(n7726), .B1(n1434), .C0(n1654), 
        .Y(N33799) );
  OAI221X2 U2412 ( .A0(n8318), .A1(n1436), .B0(n7737), .B1(n1438), .C0(n1657), 
        .Y(N33798) );
  OAI221X2 U2416 ( .A0(n8313), .A1(n1440), .B0(n7717), .B1(n1442), .C0(n1660), 
        .Y(N33797) );
  OAI221X2 U2420 ( .A0(n8313), .A1(n1444), .B0(n7717), .B1(n1446), .C0(n1663), 
        .Y(N33796) );
  OAI221X2 U2424 ( .A0(n8313), .A1(n1448), .B0(n7717), .B1(n1450), .C0(n1666), 
        .Y(N33795) );
  OAI221X2 U2428 ( .A0(n8313), .A1(n1452), .B0(n7717), .B1(n1454), .C0(n1669), 
        .Y(N33794) );
  OAI221X2 U2432 ( .A0(n8313), .A1(n1456), .B0(n7717), .B1(n1458), .C0(n1672), 
        .Y(N33793) );
  OAI221X2 U2436 ( .A0(n8313), .A1(n1460), .B0(n7717), .B1(n1462), .C0(n1675), 
        .Y(N33792) );
  OAI221X2 U2440 ( .A0(n8313), .A1(n1464), .B0(n7717), .B1(n1466), .C0(n1678), 
        .Y(N33791) );
  OAI221X2 U2444 ( .A0(n8313), .A1(n1468), .B0(n7717), .B1(n1470), .C0(n1681), 
        .Y(N33790) );
  OAI221X2 U2448 ( .A0(n8313), .A1(n1472), .B0(n7717), .B1(n1474), .C0(n1684), 
        .Y(N33789) );
  OAI221X2 U2452 ( .A0(n8313), .A1(n1476), .B0(n7717), .B1(n1478), .C0(n1687), 
        .Y(N33788) );
  OAI221X2 U2456 ( .A0(n8313), .A1(n1480), .B0(n7717), .B1(n1482), .C0(n1690), 
        .Y(N33787) );
  OAI221X2 U2460 ( .A0(n8313), .A1(n1484), .B0(n7717), .B1(n1486), .C0(n1693), 
        .Y(N33786) );
  OAI221X2 U2464 ( .A0(n8313), .A1(n1488), .B0(n7717), .B1(n1490), .C0(n1696), 
        .Y(N33785) );
  OAI221X2 U2468 ( .A0(n8314), .A1(n1492), .B0(n7718), .B1(n1494), .C0(n1699), 
        .Y(N33784) );
  OAI221X2 U2472 ( .A0(n8314), .A1(n1496), .B0(n7718), .B1(n1498), .C0(n1702), 
        .Y(N33783) );
  OAI221X2 U2476 ( .A0(n8314), .A1(n1500), .B0(n7718), .B1(n1502), .C0(n1705), 
        .Y(N33782) );
  OAI221X2 U2480 ( .A0(n8314), .A1(n1504), .B0(n7718), .B1(n1506), .C0(n1708), 
        .Y(N33781) );
  OAI221X2 U2484 ( .A0(n8314), .A1(n1508), .B0(n7718), .B1(n1510), .C0(n1711), 
        .Y(N33780) );
  OAI221X2 U2488 ( .A0(n8314), .A1(n1512), .B0(n7718), .B1(n1514), .C0(n1714), 
        .Y(N33779) );
  OAI221X2 U2492 ( .A0(n8314), .A1(n1516), .B0(n7718), .B1(n1518), .C0(n1717), 
        .Y(N33778) );
  OAI221X2 U2496 ( .A0(n8314), .A1(n1520), .B0(n7718), .B1(n1522), .C0(n1720), 
        .Y(N33777) );
  OAI221X2 U2500 ( .A0(n8314), .A1(n1524), .B0(n7718), .B1(n1526), .C0(n1723), 
        .Y(N33776) );
  OAI221X2 U2504 ( .A0(n8314), .A1(n1528), .B0(n7718), .B1(n1530), .C0(n1726), 
        .Y(N33775) );
  OAI221X2 U2508 ( .A0(n8314), .A1(n1532), .B0(n7718), .B1(n1534), .C0(n1729), 
        .Y(N33774) );
  OAI211X2 U2528 ( .A0(n7751), .A1(n1296), .B0(n1744), .C0(n1745), .Y(N33769)
         );
  OAI211X2 U2538 ( .A0(n7751), .A1(n1300), .B0(n1757), .C0(n1758), .Y(N33768)
         );
  OAI211X2 U3148 ( .A0(n7752), .A1(n1544), .B0(n2306), .C0(n2307), .Y(N33707)
         );
  GSIM_DW01_inc_0 add_272 ( .A(outCount), .SUM({N35115, N35114, N35113, N35112, 
        N35111, N35110, N35109, N35108, N35107, N35106, N35105, N35104, N35103, 
        N35102, N35101, N35100, N35099, N35098, N35097, N35096, N35095, N35094, 
        N35093, N35092, N35091, N35090, N35089, N35088, N35087, N35086, N35085, 
        N35084}) );
  GSIM_DW01_inc_1 add_258 ( .A(iCount), .SUM({N35048, N35047, N35046, N35045, 
        N35044, N35043, N35042, N35041, N35040, N35039, N35038, N35037, N35036, 
        N35035, N35034, N35033, N35032, N35031, N35030, N35029, N35028, N35027, 
        N35026, N35025, N35024, N35023, N35022, N35021, N35020, N35019, N35018, 
        N35017}) );
  GSIM_DW_div_tc_0 div_194 ( .a({N34729, N34728, N34727, N34726, N34725, 
        N34724, N34723, N34722, N34721, N34720, N34719, N34718, N34717, N34716, 
        N34715, N34714, N34713, N34712, N34711, N34710, N34709, N34708, N34707, 
        N34706, N34705, N34704, N34703, N34702, N34701, N34700, N34699, N34698, 
        N34697, N34696, N34695, N34694, N34693, N34692, N34691, N34690, N34689, 
        N34688, N34687, N34686, N34685, N34684, N34683, N34682, N34681, N34680, 
        N34679, N34678, N34677, N34676, N34675, N34674, N34673, N34672, N34671, 
        N34670, N34669, N34668, N34667, N34666}), .b({1'b0, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b0}), .quotient({N34793, N34792, N34791, N34790, N34789, 
        N34788, N34787, N34786, N34785, N34784, N34783, N34782, N34781, N34780, 
        N34779, N34778, N34777, N34776, N34775, N34774, N34773, N34772, N34771, 
        N34770, N34769, N34768, N34767, N34766, N34765, N34764, N34763, N34762, 
        N34761, N34760, N34759, N34758, N34757, N34756, N34755, N34754, N34753, 
        N34752, N34751, N34750, N34749, N34748, N34747, N34746, N34745, N34744, 
        N34743, N34742, N34741, N34740, N34739, N34738, N34737, N34736, N34735, 
        N34734, N34733, N34732, N34731, N34730}) );
  GSIM_DW_div_tc_1 div_191 ( .a({N33641, N33640, N33639, N33638, N33637, 
        N33636, N33635, N33634, N33633, N33632, N33631, N33630, N33629, N33628, 
        N33627, N33626, N33625, N33624, N33623, N33622, N33621, N33620, N33619, 
        N33618, N33617, N33616, N33615, N33614, N33613, N33612, N33611, N33610, 
        N33609, N33608, N33607, N33606, N33605, N33604, N33603, N33602, N33601, 
        N33600, N33599, N33598, N33597, N33596, N33595, N33594, N33593, N33592, 
        N33591, N33590, N33589, N33588, N33587, N33586, N33585, N33584, N33583, 
        N33582, N33581, N33580, N33579, N33578}), .b({1'b0, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b0}), .quotient({N33705, N33704, N33703, N33702, N33701, 
        N33700, N33699, N33698, N33697, N33696, N33695, N33694, N33693, N33692, 
        N33691, N33690, N33689, N33688, N33687, N33686, N33685, N33684, N33683, 
        N33682, N33681, N33680, N33679, N33678, N33677, N33676, N33675, N33674, 
        N33673, N33672, N33671, N33670, N33669, N33668, N33667, N33666, N33665, 
        N33664, N33663, N33662, N33661, N33660, N33659, N33658, N33657, N33656, 
        N33655, N33654, N33653, N33652, N33651, N33650, N33649, N33648, N33647, 
        N33646, N33645, N33644, N33643, N33642}) );
  GSIM_DW_div_tc_2 div_188 ( .a({N32681, N32680, N32679, N32678, N32677, 
        N32676, N32675, N32674, N32673, N32672, N32671, N32670, N32669, N32668, 
        N32667, N32666, N32665, N32664, N32663, N32662, N32661, N32660, N32659, 
        N32658, N32657, N32656, N32655, N32654, N32653, N32652, N32651, N32650, 
        N32649, N32648, N32647, N32646, N32645, N32644, N32643, N32642, N32641, 
        N32640, N32639, N32638, N32637, N32636, N32635, N32634, N32633, N32632, 
        N32631, N32630, N32629, N32628, N32627, N32626, N32625, N32624, N32623, 
        N32622, N32621, N32620, N32619, N32618}), .b({1'b0, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b0}), .quotient({N32745, N32744, N32743, N32742, N32741, 
        N32740, N32739, N32738, N32737, N32736, N32735, N32734, N32733, N32732, 
        N32731, N32730, N32729, N32728, N32727, N32726, N32725, N32724, N32723, 
        N32722, N32721, N32720, N32719, N32718, N32717, N32716, N32715, N32714, 
        N32713, N32712, N32711, N32710, N32709, N32708, N32707, N32706, N32705, 
        N32704, N32703, N32702, N32701, N32700, N32699, N32698, N32697, N32696, 
        N32695, N32694, N32693, N32692, N32691, N32690, N32689, N32688, N32687, 
        N32686, N32685, N32684, N32683, N32682}) );
  GSIM_DW_div_tc_3 div_185 ( .a({N31913, N31912, N31911, N31910, N31909, 
        N31908, N31907, N31906, N31905, N31904, N31903, N31902, N31901, N31900, 
        N31899, N31898, N31897, N31896, N31895, N31894, N31893, N31892, N31891, 
        N31890, N31889, N31888, N31887, N31886, N31885, N31884, N31883, N31882, 
        N31881, N31880, N31879, N31878, N31877, N31876, N31875, N31874, N31873, 
        N31872, N31871, N31870, N31869, N31868, N31867, N31866, N31865, N31864, 
        N31863, N31862, N31861, N31860, N31859, N31858, N31857, N31856, N31855, 
        N31854, N31853, N31852, N31851, N31850}), .b({1'b0, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b0}), .quotient({N31977, N31976, N31975, N31974, N31973, 
        N31972, N31971, N31970, N31969, N31968, N31967, N31966, N31965, N31964, 
        N31963, N31962, N31961, N31960, N31959, N31958, N31957, N31956, N31955, 
        N31954, N31953, N31952, N31951, N31950, N31949, N31948, N31947, N31946, 
        N31945, N31944, N31943, N31942, N31941, N31940, N31939, N31938, N31937, 
        N31936, N31935, N31934, N31933, N31932, N31931, N31930, N31929, N31928, 
        N31927, N31926, N31925, N31924, N31923, N31922, N31921, N31920, N31919, 
        N31918, N31917, N31916, N31915, N31914}) );
  GSIM_DW_div_tc_4 div_182 ( .a({N31337, N31336, N31335, N31334, N31333, 
        N31332, N31331, N31330, N31329, N31328, N31327, N31326, N31325, N31324, 
        N31323, N31322, N31321, N31320, N31319, N31318, N31317, N31316, N31315, 
        N31314, N31313, N31312, N31311, N31310, N31309, N31308, N31307, N31306, 
        N31305, N31304, N31303, N31302, N31301, N31300, N31299, N31298, N31297, 
        N31296, N31295, N31294, N31293, N31292, N31291, N31290, N31289, N31288, 
        N31287, N31286, N31285, N31284, N31283, N31282, N31281, N31280, N31279, 
        N31278, N31277, N31276, N31275, N31274}), .b({1'b0, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b0}), .quotient({N31401, N31400, N31399, N31398, N31397, 
        N31396, N31395, N31394, N31393, N31392, N31391, N31390, N31389, N31388, 
        N31387, N31386, N31385, N31384, N31383, N31382, N31381, N31380, N31379, 
        N31378, N31377, N31376, N31375, N31374, N31373, N31372, N31371, N31370, 
        N31369, N31368, N31367, N31366, N31365, N31364, N31363, N31362, N31361, 
        N31360, N31359, N31358, N31357, N31356, N31355, N31354, N31353, N31352, 
        N31351, N31350, N31349, N31348, N31347, N31346, N31345, N31344, N31343, 
        N31342, N31341, N31340, N31339, N31338}) );
  GSIM_DW_div_tc_5 div_179 ( .a({N30377, N30376, N30375, N30374, N30373, 
        N30372, N30371, N30370, N30369, N30368, N30367, N30366, N30365, N30364, 
        N30363, N30362, N30361, N30360, N30359, N30358, N30357, N30356, N30355, 
        N30354, N30353, N30352, N30351, N30350, N30349, N30348, N30347, N30346, 
        N30345, N30344, N30343, N30342, N30341, N30340, N30339, N30338, N30337, 
        N30336, N30335, N30334, N30333, N30332, N30331, N30330, N30329, N30328, 
        N30327, N30326, N30325, N30324, N30323, N30322, N30321, N30320, N30319, 
        N30318, N30317, N30316, N30315, N30314}), .b({1'b0, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b0}), .quotient({N30441, N30440, N30439, N30438, N30437, 
        N30436, N30435, N30434, N30433, N30432, N30431, N30430, N30429, N30428, 
        N30427, N30426, N30425, N30424, N30423, N30422, N30421, N30420, N30419, 
        N30418, N30417, N30416, N30415, N30414, N30413, N30412, N30411, N30410, 
        N30409, N30408, N30407, N30406, N30405, N30404, N30403, N30402, N30401, 
        N30400, N30399, N30398, N30397, N30396, N30395, N30394, N30393, N30392, 
        N30391, N30390, N30389, N30388, N30387, N30386, N30385, N30384, N30383, 
        N30382, N30381, N30380, N30379, N30378}) );
  GSIM_DW_div_tc_6 div_176 ( .a({N29609, N29608, N29607, N29606, N29605, 
        N29604, N29603, N29602, N29601, N29600, N29599, N29598, N29597, N29596, 
        N29595, N29594, N29593, N29592, N29591, N29590, N29589, N29588, N29587, 
        N29586, N29585, N29584, N29583, N29582, N29581, N29580, N29579, N29578, 
        N29577, N29576, N29575, N29574, N29573, N29572, N29571, N29570, N29569, 
        N29568, N29567, N29566, N29565, N29564, N29563, N29562, N29561, N29560, 
        N29559, N29558, N29557, N29556, N29555, N29554, N29553, N29552, N29551, 
        N29550, N29549, N29548, N29547, N29546}), .b({1'b0, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b0}), .quotient({N29673, N29672, N29671, N29670, N29669, 
        N29668, N29667, N29666, N29665, N29664, N29663, N29662, N29661, N29660, 
        N29659, N29658, N29657, N29656, N29655, N29654, N29653, N29652, N29651, 
        N29650, N29649, N29648, N29647, N29646, N29645, N29644, N29643, N29642, 
        N29641, N29640, N29639, N29638, N29637, N29636, N29635, N29634, N29633, 
        N29632, N29631, N29630, N29629, N29628, N29627, N29626, N29625, N29624, 
        N29623, N29622, N29621, N29620, N29619, N29618, N29617, N29616, N29615, 
        N29614, N29613, N29612, N29611, N29610}) );
  GSIM_DW_div_tc_7 div_163 ( .a({N25537, N25538, N25539, N25540, N25541, 
        N25542, N25543, N25544, N25545, N25546, N25547, N25548, N25549, N25550, 
        N25551, N25552, N25553, N25554, N25555, N25556, N25557, N25558, N25559, 
        N25560, N25561, N25562, N25563, N25564, N25565, N25566, N25567, N25568, 
        N25569, N25570, N25571, N25572, N25573, N25574, N25575, N25576, N25577, 
        N25578, N25579, N25580, N25581, N25582, N25583, N25584, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .b({1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0}), .quotient({
        N25664, SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, N25661, 
        N25660, N25659, N25658, N25657, N25656, N25655, N25654, N25653, N25652, 
        N25651, N25650, N25649, N25648, N25647, N25646, N25645, N25644, N25643, 
        N25642, N25641, N25640, N25639, N25638, N25637, N25636, N25635, N25634, 
        N25633, N25632, N25631, N25630, N25629, N25628, N25627, N25626, N25625, 
        N25624, N25623, N25622, N25621, N25620, N25619, N25618, N25617, N25616, 
        N25615, N25614, N25613, N25612, N25611, N25610, N25609, N25608, N25607, 
        N25606, N25605, N25604, N25603, N25602, N25601}) );
  GSIM_DW01_inc_10 add_104 ( .A({inCount[31:4], n8411, n8412, n8413, n8414}), 
        .SUM({N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, 
        N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, 
        N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, 
        N1775, N1774, N1773}) );
  GSIM_DW01_inc_11 r1198 ( .A({xCount[31:4], n8407, n8408, n8409, n8410}), 
        .SUM({N34908, N34907, N34906, N34905, N34904, N34903, N34902, N34901, 
        N34900, N34899, N34898, N34897, N34896, N34895, N34894, N34893, N34892, 
        N34891, N34890, N34889, N34888, N34887, N34886, N34885, N34884, N34883, 
        N34882, N34881, N34880, N34879, N34878, N34877}) );
  GSIM_DW_mult_tc_21 mult_194_3 ( .a({1'b0, 1'b1, 1'b1, 1'b0, 1'b1}), .b({
        N33897, N33896, N33895, N33894, N33893, N33892, N33891, N33890, N33889, 
        N33888, N33887, N33886, N33885, N33884, N33883, N33882, N33881, N33880, 
        N33879, N33878, N33877, N33876, N33875, N33874, N33873, N33872, N33871, 
        N33870, N33869, N33868, N33867, N33866, N33865, N33864, N33863, N33862, 
        N33861, N33860, N33859, N33858, N33857, N33856, N33855, N33854, N33853, 
        N33852, N33851, N33850, N33849, N33848, N33847, N33846, N33845, N33844, 
        N33843, N33842, N33841, N33840, N33839, N33838, N33837, N33836, N33835, 
        N33834}), .product({SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, N34345, N34344, N34343, N34342, N34341, 
        N34340, N34339, N34338, N34337, N34336, N34335, N34334, N34333, N34332, 
        N34331, N34330, N34329, N34328, N34327, N34326, N34325, N34324, N34323, 
        N34322, N34321, N34320, N34319, N34318, N34317, N34316, N34315, N34314, 
        N34313, N34312, N34311, N34310, N34309, N34308, N34307, N34306, N34305, 
        N34304, N34303, N34302, N34301, N34300, N34299, N34298, N34297, N34296, 
        N34295, N34294, N34293, N34292, N34291, N34290, N34289, N34288, N34287, 
        N34286, N34285, N34284, N34283, N34282}) );
  GSIM_DW_mult_tc_20 mult_194_5 ( .a({1'b1, 1'b0, 1'b1, 1'b0}), .b({N34025, 
        N34024, N34023, N34022, N34021, N34020, N34019, N34018, N34017, N34016, 
        N34015, N34014, N34013, N34012, N34011, N34010, N34009, N34008, N34007, 
        N34006, N34005, N34004, N34003, N34002, N34001, N34000, N33999, N33998, 
        N33997, N33996, N33995, N33994, N33993, N33992, N33991, N33990, N33989, 
        N33988, N33987, N33986, N33985, N33984, N33983, N33982, N33981, N33980, 
        N33979, N33978, N33977, N33976, N33975, N33974, N33973, N33972, N33971, 
        N33970, N33969, N33968, N33967, N33966, N33965, N33964, N33963, N33962}), .product({SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, N34601, N34600, 
        N34599, N34598, N34597, N34596, N34595, N34594, N34593, N34592, N34591, 
        N34590, N34589, N34588, N34587, N34586, N34585, N34584, N34583, N34582, 
        N34581, N34580, N34579, N34578, N34577, N34576, N34575, N34574, N34573, 
        N34572, N34571, N34570, N34569, N34568, N34567, N34566, N34565, N34564, 
        N34563, N34562, N34561, N34560, N34559, N34558, N34557, N34556, N34555, 
        N34554, N34553, N34552, N34551, N34550, N34549, N34548, N34547, N34546, 
        N34545, N34544, N34543, N34542, N34541, N34540, N34539, 
        SYNOPSYS_UNCONNECTED__11}) );
  GSIM_DW_mult_tc_19 mult_194_2 ( .a({1'b1, 1'b0, 1'b1, 1'b0}), .b({N33833, 
        N33832, N33831, N33830, N33829, N33828, N33827, N33826, N33825, N33824, 
        N33823, N33822, N33821, N33820, N33819, N33818, N33817, N33816, N33815, 
        N33814, N33813, N33812, N33811, N33810, N33809, N33808, N33807, N33806, 
        N33805, N33804, N33803, N33802, N33801, N33800, N33799, N33798, N33797, 
        N33796, N33795, N33794, N33793, N33792, N33791, N33790, N33789, N33788, 
        N33787, N33786, N33785, N33784, N33783, N33782, N33781, N33780, N33779, 
        N33778, N33777, N33776, N33775, N33774, N33773, N33772, N33771, N33770}), .product({SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, N34217, N34216, 
        N34215, N34214, N34213, N34212, N34211, N34210, N34209, N34208, N34207, 
        N34206, N34205, N34204, N34203, N34202, N34201, N34200, N34199, N34198, 
        N34197, N34196, N34195, N34194, N34193, N34192, N34191, N34190, N34189, 
        N34188, N34187, N34186, N34185, N34184, N34183, N34182, N34181, N34180, 
        N34179, N34178, N34177, N34176, N34175, N34174, N34173, N34172, N34171, 
        N34170, N34169, N34168, N34167, N34166, N34165, N34164, N34163, N34162, 
        N34161, N34160, N34159, N34158, N34157, N34156, N34155, 
        SYNOPSYS_UNCONNECTED__16}) );
  GSIM_DW01_add_501 add_5_root_add_0_root_add_194_9 ( .A({N28833, N28834, 
        N28835, N28836, N28837, N28838, N28839, N28840, N28841, N28842, N28843, 
        N28844, N28845, N28846, N28847, N28848, N28849, N28850, N28851, N28852, 
        N28853, N28854, N28855, N28856, N28857, N28858, N28859, N28860, N28861, 
        N28862, N28863, N28864, N28865, N28866, N28867, N28868, N28869, N28870, 
        N28871, N28872, N28873, N28874, N28875, N28876, N28877, N28878, N28879, 
        N28880, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N34217, N34216, N34215, 
        N34214, N34213, N34212, N34211, N34210, N34209, N34208, N34207, N34206, 
        N34205, N34204, N34203, N34202, N34201, N34200, N34199, N34198, N34197, 
        N34196, N34195, N34194, N34193, N34192, N34191, N34190, N34189, N34188, 
        N34187, N34186, N34185, N34184, N34183, N34182, N34181, N34180, N34179, 
        N34178, N34177, N34176, N34175, N34174, N34173, N34172, N34171, N34170, 
        N34169, N34168, N34167, N34166, N34165, N34164, N34163, N34162, N34161, 
        N34160, N34159, N34158, N34157, N34156, N34155, 1'b0}), .CI(1'b0), 
        .SUM({N34409, N34408, N34407, N34406, N34405, N34404, N34403, N34402, 
        N34401, N34400, N34399, N34398, N34397, N34396, N34395, N34394, N34393, 
        N34392, N34391, N34390, N34389, N34388, N34387, N34386, N34385, N34384, 
        N34383, N34382, N34381, N34380, N34379, N34378, N34377, N34376, N34375, 
        N34374, N34373, N34372, N34371, N34370, N34369, N34368, N34367, N34366, 
        N34365, N34364, N34363, N34362, N34361, N34360, N34359, N34358, N34357, 
        N34356, N34355, N34354, N34353, N34352, N34351, N34350, N34349, N34348, 
        N34347, SYNOPSYS_UNCONNECTED__17}) );
  GSIM_DW01_add_500 add_4_root_add_0_root_add_194_9 ( .A({N34601, N34600, 
        N34599, N34598, N34597, N34596, N34595, N34594, N34593, N34592, N34591, 
        N34590, N34589, N34588, N34587, N34586, N34585, N34584, N34583, N34582, 
        N34581, N34580, N34579, N34578, N34577, N34576, N34575, N34574, N34573, 
        N34572, N34571, N34570, N34569, N34568, N34567, N34566, N34565, N34564, 
        N34563, N34562, N34561, N34560, N34559, N34558, N34557, N34556, N34555, 
        N34554, N34553, N34552, N34551, N34550, N34549, N34548, N34547, N34546, 
        N34545, N34544, N34543, N34542, N34541, N34540, N34539, 1'b0}), .B({
        N34409, N34408, N34407, N34406, N34405, N34404, N34403, N34402, N34401, 
        N34400, N34399, N34398, N34397, N34396, N34395, N34394, N34393, N34392, 
        N34391, N34390, N34389, N34388, N34387, N34386, N34385, N34384, N34383, 
        N34382, N34381, N34380, N34379, N34378, N34377, N34376, N34375, N34374, 
        N34373, N34372, N34371, N34370, N34369, N34368, N34367, N34366, N34365, 
        N34364, N34363, N34362, N34361, N34360, N34359, N34358, N34357, N34356, 
        N34355, N34354, N34353, N34352, N34351, N34350, N34349, N34348, N34347, 
        1'b0}), .CI(1'b0), .SUM({N34281, N34280, N34279, N34278, N34277, 
        N34276, N34275, N34274, N34273, N34272, N34271, N34270, N34269, N34268, 
        N34267, N34266, N34265, N34264, N34263, N34262, N34261, N34260, N34259, 
        N34258, N34257, N34256, N34255, N34254, N34253, N34252, N34251, N34250, 
        N34249, N34248, N34247, N34246, N34245, N34244, N34243, N34242, N34241, 
        N34240, N34239, N34238, N34237, N34236, N34235, N34234, N34233, N34232, 
        N34231, N34230, N34229, N34228, N34227, N34226, N34225, N34224, N34223, 
        N34222, N34221, N34220, N34219, SYNOPSYS_UNCONNECTED__18}) );
  GSIM_DW_mult_tc_18 mult_194_4 ( .a({1'b0, 1'b1, 1'b1, 1'b0, 1'b1}), .b({
        N33961, N33960, N33959, N33958, N33957, N33956, N33955, N33954, N33953, 
        N33952, N33951, N33950, N33949, N33948, N33947, N33946, N33945, N33944, 
        N33943, N33942, N33941, N33940, N33939, N33938, N33937, N33936, N33935, 
        N33934, N33933, N33932, N33931, N33930, N33929, N33928, N33927, N33926, 
        N33925, N33924, N33923, N33922, N33921, N33920, N33919, N33918, N33917, 
        N33916, N33915, N33914, N33913, N33912, N33911, N33910, N33909, N33908, 
        N33907, N33906, N33905, N33904, N33903, N33902, N33901, N33900, N33899, 
        N33898}), .product({SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, N34473, N34472, N34471, N34470, N34469, 
        N34468, N34467, N34466, N34465, N34464, N34463, N34462, N34461, N34460, 
        N34459, N34458, N34457, N34456, N34455, N34454, N34453, N34452, N34451, 
        N34450, N34449, N34448, N34447, N34446, N34445, N34444, N34443, N34442, 
        N34441, N34440, N34439, N34438, N34437, N34436, N34435, N34434, N34433, 
        N34432, N34431, N34430, N34429, N34428, N34427, N34426, N34425, N34424, 
        N34423, N34422, N34421, N34420, N34419, N34418, N34417, N34416, N34415, 
        N34414, N34413, N34412, N34411, N34410}) );
  GSIM_DW01_add_499 add_3_root_add_0_root_add_194_9 ( .A({N34281, N34280, 
        N34279, N34278, N34277, N34276, N34275, N34274, N34273, N34272, N34271, 
        N34270, N34269, N34268, N34267, N34266, N34265, N34264, N34263, N34262, 
        N34261, N34260, N34259, N34258, N34257, N34256, N34255, N34254, N34253, 
        N34252, N34251, N34250, N34249, N34248, N34247, N34246, N34245, N34244, 
        N34243, N34242, N34241, N34240, N34239, N34238, N34237, N34236, N34235, 
        N34234, N34233, N34232, N34231, N34230, N34229, N34228, N34227, N34226, 
        N34225, N34224, N34223, N34222, N34221, N34220, N34219, 1'b0}), .B({
        N34473, N34472, N34471, N34470, N34469, N34468, N34467, N34466, N34465, 
        N34464, N34463, N34462, N34461, N34460, N34459, N34458, N34457, N34456, 
        N34455, N34454, N34453, N34452, N34451, N34450, N34449, N34448, N34447, 
        N34446, N34445, N34444, N34443, N34442, N34441, N34440, N34439, N34438, 
        N34437, N34436, N34435, N34434, N34433, N34432, N34431, N34430, N34429, 
        N34428, N34427, N34426, N34425, N34424, N34423, N34422, N34421, N34420, 
        N34419, N34418, N34417, N34416, N34415, N34414, N34413, N34412, N34411, 
        N34410}), .CI(1'b0), .SUM({N34665, N34664, N34663, N34662, N34661, 
        N34660, N34659, N34658, N34657, N34656, N34655, N34654, N34653, N34652, 
        N34651, N34650, N34649, N34648, N34647, N34646, N34645, N34644, N34643, 
        N34642, N34641, N34640, N34639, N34638, N34637, N34636, N34635, N34634, 
        N34633, N34632, N34631, N34630, N34629, N34628, N34627, N34626, N34625, 
        N34624, N34623, N34622, N34621, N34620, N34619, N34618, N34617, N34616, 
        N34615, N34614, N34613, N34612, N34611, N34610, N34609, N34608, N34607, 
        N34606, N34605, N34604, N34603, N34602}) );
  GSIM_DW01_add_498 add_2_root_add_0_root_add_194_9 ( .A({N34345, N34344, 
        N34343, N34342, N34341, N34340, N34339, N34338, N34337, N34336, N34335, 
        N34334, N34333, N34332, N34331, N34330, N34329, N34328, N34327, N34326, 
        N34325, N34324, N34323, N34322, N34321, N34320, N34319, N34318, N34317, 
        N34316, N34315, N34314, N34313, N34312, N34311, N34310, N34309, N34308, 
        N34307, N34306, N34305, N34304, N34303, N34302, N34301, N34300, N34299, 
        N34298, N34297, N34296, N34295, N34294, N34293, N34292, N34291, N34290, 
        N34289, N34288, N34287, N34286, N34285, N34284, N34283, N34282}), .B({
        N34665, N34664, N34663, N34662, N34661, N34660, N34659, N34658, N34657, 
        N34656, N34655, N34654, N34653, N34652, N34651, N34650, N34649, N34648, 
        N34647, N34646, N34645, N34644, N34643, N34642, N34641, N34640, N34639, 
        N34638, N34637, N34636, N34635, N34634, N34633, N34632, N34631, N34630, 
        N34629, N34628, N34627, N34626, N34625, N34624, N34623, N34622, N34621, 
        N34620, N34619, N34618, N34617, N34616, N34615, N34614, N34613, N34612, 
        N34611, N34610, N34609, N34608, N34607, N34606, N34605, N34604, N34603, 
        N34602}), .CI(1'b0), .SUM({N34153, N34152, N34151, N34150, N34149, 
        N34148, N34147, N34146, N34145, N34144, N34143, N34142, N34141, N34140, 
        N34139, N34138, N34137, N34136, N34135, N34134, N34133, N34132, N34131, 
        N34130, N34129, N34128, N34127, N34126, N34125, N34124, N34123, N34122, 
        N34121, N34120, N34119, N34118, N34117, N34116, N34115, N34114, N34113, 
        N34112, N34111, N34110, N34109, N34108, N34107, N34106, N34105, N34104, 
        N34103, N34102, N34101, N34100, N34099, N34098, N34097, N34096, N34095, 
        N34094, N34093, N34092, N34091, N34090}) );
  GSIM_DW01_add_497 add_1_root_add_0_root_add_194_9 ( .A({N34153, N34152, 
        N34151, N34150, N34149, N34148, N34147, N34146, N34145, N34144, N34143, 
        N34142, N34141, N34140, N34139, N34138, N34137, N34136, N34135, N34134, 
        N34133, N34132, N34131, N34130, N34129, N34128, N34127, N34126, N34125, 
        N34124, N34123, N34122, N34121, N34120, N34119, N34118, N34117, N34116, 
        N34115, N34114, N34113, N34112, N34111, N34110, N34109, N34108, N34107, 
        N34106, N34105, N34104, N34103, N34102, N34101, N34100, N34099, N34098, 
        N34097, N34096, N34095, N34094, N34093, N34092, N34091, N34090}), .B({
        N33769, N33768, N33767, N33766, N33765, N33764, N33763, N33762, N33761, 
        N33760, N33759, N33758, N33757, N33756, N33755, N33754, N33753, N33752, 
        N33751, N33750, N33749, N33748, N33747, N33746, N33745, N33744, N33743, 
        N33742, N33741, N33740, N33739, N33738, N33737, N33736, N33735, N33734, 
        N33733, N33732, N33731, N33730, N33729, N33728, N33727, N33726, N33725, 
        N33724, N33723, N33722, N33721, N33720, N33719, N33718, N33717, N33716, 
        N33715, N33714, N33713, N33712, N33711, N33710, N33709, N33708, N33707, 
        N33706}), .CI(1'b0), .SUM({N34537, N34536, N34535, N34534, N34533, 
        N34532, N34531, N34530, N34529, N34528, N34527, N34526, N34525, N34524, 
        N34523, N34522, N34521, N34520, N34519, N34518, N34517, N34516, N34515, 
        N34514, N34513, N34512, N34511, N34510, N34509, N34508, N34507, N34506, 
        N34505, N34504, N34503, N34502, N34501, N34500, N34499, N34498, N34497, 
        N34496, N34495, N34494, N34493, N34492, N34491, N34490, N34489, N34488, 
        N34487, N34486, N34485, N34484, N34483, N34482, N34481, N34480, N34479, 
        N34478, N34477, N34476, N34475, N34474}) );
  GSIM_DW01_add_496 add_0_root_add_0_root_add_194_9 ( .A({N34089, N34088, 
        N34087, N34086, N34085, N34084, N34083, N34082, N34081, N34080, N34079, 
        N34078, N34077, N34076, N34075, N34074, N34073, N34072, N34071, N34070, 
        N34069, N34068, N34067, N34066, N34065, N34064, N34063, N34062, N34061, 
        N34060, N34059, N34058, N34057, N34056, N34055, N34054, N34053, N34052, 
        N34051, N34050, N34049, N34048, N34047, N34046, N34045, N34044, N34043, 
        N34042, N34041, N34040, N34039, N34038, N34037, N34036, N34035, N34034, 
        N34033, N34032, N34031, N34030, N34029, N34028, N34027, N34026}), .B({
        N34537, N34536, N34535, N34534, N34533, N34532, N34531, N34530, N34529, 
        N34528, N34527, N34526, N34525, N34524, N34523, N34522, N34521, N34520, 
        N34519, N34518, N34517, N34516, N34515, N34514, N34513, N34512, N34511, 
        N34510, N34509, N34508, N34507, N34506, N34505, N34504, N34503, N34502, 
        N34501, N34500, N34499, N34498, N34497, N34496, N34495, N34494, N34493, 
        N34492, N34491, N34490, N34489, N34488, N34487, N34486, N34485, N34484, 
        N34483, N34482, N34481, N34480, N34479, N34478, N34477, N34476, N34475, 
        N34474}), .CI(1'b0), .SUM({N34729, N34728, N34727, N34726, N34725, 
        N34724, N34723, N34722, N34721, N34720, N34719, N34718, N34717, N34716, 
        N34715, N34714, N34713, N34712, N34711, N34710, N34709, N34708, N34707, 
        N34706, N34705, N34704, N34703, N34702, N34701, N34700, N34699, N34698, 
        N34697, N34696, N34695, N34694, N34693, N34692, N34691, N34690, N34689, 
        N34688, N34687, N34686, N34685, N34684, N34683, N34682, N34681, N34680, 
        N34679, N34678, N34677, N34676, N34675, N34674, N34673, N34672, N34671, 
        N34670, N34669, N34668, N34667, N34666}) );
  GSIM_DW_mult_tc_3 mult_182 ( .a({1'b1, 1'b0, 1'b1, 1'b0}), .b({N33833, 
        N33832, N33831, N33830, N33829, N33828, N33827, N33826, N33825, N33824, 
        N33823, N33822, N33821, N33820, N33819, N33818, N33817, N33816, N33815, 
        N33814, N33813, N33812, N33811, N33810, N33809, N33808, N33807, N33806, 
        N33805, N33804, N33803, N33802, N33801, N33800, N33799, N33798, N33797, 
        N33796, N33795, N33794, N33793, N33792, N33791, N33790, N33789, N33788, 
        N33787, N33786, N33785, N33784, N33783, N33782, N33781, N33780, N33779, 
        N33778, N33777, N33776, N33775, N33774, N33773, N33772, N33771, N33770}), .product({SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, N30825, N30824, 
        N30823, N30822, N30821, N30820, N30819, N30818, N30817, N30816, N30815, 
        N30814, N30813, N30812, N30811, N30810, N30809, N30808, N30807, N30806, 
        N30805, N30804, N30803, N30802, N30801, N30800, N30799, N30798, N30797, 
        N30796, N30795, N30794, N30793, N30792, N30791, N30790, N30789, N30788, 
        N30787, N30786, N30785, N30784, N30783, N30782, N30781, N30780, N30779, 
        N30778, N30777, N30776, N30775, N30774, N30773, N30772, N30771, N30770, 
        N30769, N30768, N30767, N30766, N30765, N30764, N30763, 
        SYNOPSYS_UNCONNECTED__28}) );
  GSIM_DW_mult_tc_2 mult_182_2 ( .a({1'b0, 1'b1, 1'b1, 1'b0, 1'b1}), .b({
        N33897, N33896, N33895, N33894, N33893, N33892, N33891, N33890, N33889, 
        N33888, N33887, N33886, N33885, N33884, N33883, N33882, N33881, N33880, 
        N33879, N33878, N33877, N33876, N33875, N33874, N33873, N33872, N33871, 
        N33870, N33869, N33868, N33867, N33866, N33865, N33864, N33863, N33862, 
        N33861, N33860, N33859, N33858, N33857, N33856, N33855, N33854, N33853, 
        N33852, N33851, N33850, N33849, N33848, N33847, N33846, N33845, N33844, 
        N33843, N33842, N33841, N33840, N33839, N33838, N33837, N33836, N33835, 
        N33834}), .product({SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, N30953, N30952, N30951, N30950, N30949, 
        N30948, N30947, N30946, N30945, N30944, N30943, N30942, N30941, N30940, 
        N30939, N30938, N30937, N30936, N30935, N30934, N30933, N30932, N30931, 
        N30930, N30929, N30928, N30927, N30926, N30925, N30924, N30923, N30922, 
        N30921, N30920, N30919, N30918, N30917, N30916, N30915, N30914, N30913, 
        N30912, N30911, N30910, N30909, N30908, N30907, N30906, N30905, N30904, 
        N30903, N30902, N30901, N30900, N30899, N30898, N30897, N30896, N30895, 
        N30894, N30893, N30892, N30891, N30890}) );
  GSIM_DW_mult_tc_1 mult_182_3 ( .a({1'b0, 1'b1, 1'b1, 1'b0, 1'b1}), .b({
        N33961, N33960, N33959, N33958, N33957, N33956, N33955, N33954, N33953, 
        N33952, N33951, N33950, N33949, N33948, N33947, N33946, N33945, N33944, 
        N33943, N33942, N33941, N33940, N33939, N33938, N33937, N33936, N33935, 
        N33934, N33933, N33932, N33931, N33930, N33929, N33928, N33927, N33926, 
        N33925, N33924, N33923, N33922, N33921, N33920, N33919, N33918, N33917, 
        N33916, N33915, N33914, N33913, N33912, N33911, N33910, N33909, N33908, 
        N33907, N33906, N33905, N33904, N33903, N33902, N33901, N33900, N33899, 
        N33898}), .product({SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, N31081, N31080, N31079, N31078, N31077, 
        N31076, N31075, N31074, N31073, N31072, N31071, N31070, N31069, N31068, 
        N31067, N31066, N31065, N31064, N31063, N31062, N31061, N31060, N31059, 
        N31058, N31057, N31056, N31055, N31054, N31053, N31052, N31051, N31050, 
        N31049, N31048, N31047, N31046, N31045, N31044, N31043, N31042, N31041, 
        N31040, N31039, N31038, N31037, N31036, N31035, N31034, N31033, N31032, 
        N31031, N31030, N31029, N31028, N31027, N31026, N31025, N31024, N31023, 
        N31022, N31021, N31020, N31019, N31018}) );
  GSIM_DW_mult_tc_0 mult_182_4 ( .a({1'b1, 1'b0, 1'b1, 1'b0}), .b({N34025, 
        N34024, N34023, N34022, N34021, N34020, N34019, N34018, N34017, N34016, 
        N34015, N34014, N34013, N34012, N34011, N34010, N34009, N34008, N34007, 
        N34006, N34005, N34004, N34003, N34002, N34001, N34000, N33999, N33998, 
        N33997, N33996, N33995, N33994, N33993, N33992, N33991, N33990, N33989, 
        N33988, N33987, N33986, N33985, N33984, N33983, N33982, N33981, N33980, 
        N33979, N33978, N33977, N33976, N33975, N33974, N33973, N33972, N33971, 
        N33970, N33969, N33968, N33967, N33966, N33965, N33964, N33963, N33962}), .product({SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, N31209, N31208, 
        N31207, N31206, N31205, N31204, N31203, N31202, N31201, N31200, N31199, 
        N31198, N31197, N31196, N31195, N31194, N31193, N31192, N31191, N31190, 
        N31189, N31188, N31187, N31186, N31185, N31184, N31183, N31182, N31181, 
        N31180, N31179, N31178, N31177, N31176, N31175, N31174, N31173, N31172, 
        N31171, N31170, N31169, N31168, N31167, N31166, N31165, N31164, N31163, 
        N31162, N31161, N31160, N31159, N31158, N31157, N31156, N31155, N31154, 
        N31153, N31152, N31151, N31150, N31149, N31148, N31147, 
        SYNOPSYS_UNCONNECTED__43}) );
  GSIM_DW01_add_476 add_3_root_add_0_root_add_182_8 ( .A({N30825, N30824, 
        N30823, N30822, N30821, N30820, N30819, N30818, N30817, N30816, N30815, 
        N30814, N30813, N30812, N30811, N30810, N30809, N30808, N30807, N30806, 
        N30805, N30804, N30803, N30802, N30801, N30800, N30799, N30798, N30797, 
        N30796, N30795, N30794, N30793, N30792, N30791, N30790, N30789, N30788, 
        N30787, N30786, N30785, N30784, N30783, N30782, N30781, N30780, N30779, 
        N30778, N30777, N30776, N30775, N30774, N30773, N30772, N30771, N30770, 
        N30769, N30768, N30767, N30766, N30765, N30764, N30763, 1'b0}), .B({
        N30953, N30952, N30951, N30950, N30949, N30948, N30947, N30946, N30945, 
        N30944, N30943, N30942, N30941, N30940, N30939, N30938, N30937, N30936, 
        N30935, N30934, N30933, N30932, N30931, N30930, N30929, N30928, N30927, 
        N30926, N30925, N30924, N30923, N30922, N30921, N30920, N30919, N30918, 
        N30917, N30916, N30915, N30914, N30913, N30912, N30911, N30910, N30909, 
        N30908, N30907, N30906, N30905, N30904, N30903, N30902, N30901, N30900, 
        N30899, N30898, N30897, N30896, N30895, N30894, N30893, N30892, N30891, 
        N30890}), .CI(1'b0), .SUM({N30889, N30888, N30887, N30886, N30885, 
        N30884, N30883, N30882, N30881, N30880, N30879, N30878, N30877, N30876, 
        N30875, N30874, N30873, N30872, N30871, N30870, N30869, N30868, N30867, 
        N30866, N30865, N30864, N30863, N30862, N30861, N30860, N30859, N30858, 
        N30857, N30856, N30855, N30854, N30853, N30852, N30851, N30850, N30849, 
        N30848, N30847, N30846, N30845, N30844, N30843, N30842, N30841, N30840, 
        N30839, N30838, N30837, N30836, N30835, N30834, N30833, N30832, N30831, 
        N30830, N30829, N30828, N30827, N30826}) );
  GSIM_DW01_add_475 add_4_root_add_0_root_add_182_8 ( .A({N28833, N28834, 
        N28835, N28836, N28837, N28838, N28839, N28840, N28841, N28842, N28843, 
        N28844, N28845, N28846, N28847, N28848, N28849, N28850, N28851, N28852, 
        N28853, N28854, N28855, N28856, N28857, N28858, N28859, N28860, N28861, 
        N28862, N28863, N28864, N28865, N28866, N28867, N28868, N28869, N28870, 
        N28871, N28872, N28873, N28874, N28875, N28876, N28877, N28878, N28879, 
        N28880, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N31209, N31208, N31207, 
        N31206, N31205, N31204, N31203, N31202, N31201, N31200, N31199, N31198, 
        N31197, N31196, N31195, N31194, N31193, N31192, N31191, N31190, N31189, 
        N31188, N31187, N31186, N31185, N31184, N31183, N31182, N31181, N31180, 
        N31179, N31178, N31177, N31176, N31175, N31174, N31173, N31172, N31171, 
        N31170, N31169, N31168, N31167, N31166, N31165, N31164, N31163, N31162, 
        N31161, N31160, N31159, N31158, N31157, N31156, N31155, N31154, N31153, 
        N31152, N31151, N31150, N31149, N31148, N31147, 1'b0}), .CI(1'b0), 
        .SUM({N31017, N31016, N31015, N31014, N31013, N31012, N31011, N31010, 
        N31009, N31008, N31007, N31006, N31005, N31004, N31003, N31002, N31001, 
        N31000, N30999, N30998, N30997, N30996, N30995, N30994, N30993, N30992, 
        N30991, N30990, N30989, N30988, N30987, N30986, N30985, N30984, N30983, 
        N30982, N30981, N30980, N30979, N30978, N30977, N30976, N30975, N30974, 
        N30973, N30972, N30971, N30970, N30969, N30968, N30967, N30966, N30965, 
        N30964, N30963, N30962, N30961, N30960, N30959, N30958, N30957, N30956, 
        N30955, SYNOPSYS_UNCONNECTED__44}) );
  GSIM_DW01_add_474 add_2_root_add_0_root_add_182_8 ( .A({N31081, N31080, 
        N31079, N31078, N31077, N31076, N31075, N31074, N31073, N31072, N31071, 
        N31070, N31069, N31068, N31067, N31066, N31065, N31064, N31063, N31062, 
        N31061, N31060, N31059, N31058, N31057, N31056, N31055, N31054, N31053, 
        N31052, N31051, N31050, N31049, N31048, N31047, N31046, N31045, N31044, 
        N31043, N31042, N31041, N31040, N31039, N31038, N31037, N31036, N31035, 
        N31034, N31033, N31032, N31031, N31030, N31029, N31028, N31027, N31026, 
        N31025, N31024, N31023, N31022, N31021, N31020, N31019, N31018}), .B({
        N31017, N31016, N31015, N31014, N31013, N31012, N31011, N31010, N31009, 
        N31008, N31007, N31006, N31005, N31004, N31003, N31002, N31001, N31000, 
        N30999, N30998, N30997, N30996, N30995, N30994, N30993, N30992, N30991, 
        N30990, N30989, N30988, N30987, N30986, N30985, N30984, N30983, N30982, 
        N30981, N30980, N30979, N30978, N30977, N30976, N30975, N30974, N30973, 
        N30972, N30971, N30970, N30969, N30968, N30967, N30966, N30965, N30964, 
        N30963, N30962, N30961, N30960, N30959, N30958, N30957, N30956, N30955, 
        1'b0}), .CI(1'b0), .SUM({N31273, N31272, N31271, N31270, N31269, 
        N31268, N31267, N31266, N31265, N31264, N31263, N31262, N31261, N31260, 
        N31259, N31258, N31257, N31256, N31255, N31254, N31253, N31252, N31251, 
        N31250, N31249, N31248, N31247, N31246, N31245, N31244, N31243, N31242, 
        N31241, N31240, N31239, N31238, N31237, N31236, N31235, N31234, N31233, 
        N31232, N31231, N31230, N31229, N31228, N31227, N31226, N31225, N31224, 
        N31223, N31222, N31221, N31220, N31219, N31218, N31217, N31216, N31215, 
        N31214, N31213, N31212, N31211, N31210}) );
  GSIM_DW01_add_473 add_1_root_add_0_root_add_182_8 ( .A({N31273, N31272, 
        N31271, N31270, N31269, N31268, N31267, N31266, N31265, N31264, N31263, 
        N31262, N31261, N31260, N31259, N31258, N31257, N31256, N31255, N31254, 
        N31253, N31252, N31251, N31250, N31249, N31248, N31247, N31246, N31245, 
        N31244, N31243, N31242, N31241, N31240, N31239, N31238, N31237, N31236, 
        N31235, N31234, N31233, N31232, N31231, N31230, N31229, N31228, N31227, 
        N31226, N31225, N31224, N31223, N31222, N31221, N31220, N31219, N31218, 
        N31217, N31216, N31215, N31214, N31213, N31212, N31211, N31210}), .B({
        N30889, N30888, N30887, N30886, N30885, N30884, N30883, N30882, N30881, 
        N30880, N30879, N30878, N30877, N30876, N30875, N30874, N30873, N30872, 
        N30871, N30870, N30869, N30868, N30867, N30866, N30865, N30864, N30863, 
        N30862, N30861, N30860, N30859, N30858, N30857, N30856, N30855, N30854, 
        N30853, N30852, N30851, N30850, N30849, N30848, N30847, N30846, N30845, 
        N30844, N30843, N30842, N30841, N30840, N30839, N30838, N30837, N30836, 
        N30835, N30834, N30833, N30832, N30831, N30830, N30829, N30828, N30827, 
        N30826}), .CI(1'b0), .SUM({N31145, N31144, N31143, N31142, N31141, 
        N31140, N31139, N31138, N31137, N31136, N31135, N31134, N31133, N31132, 
        N31131, N31130, N31129, N31128, N31127, N31126, N31125, N31124, N31123, 
        N31122, N31121, N31120, N31119, N31118, N31117, N31116, N31115, N31114, 
        N31113, N31112, N31111, N31110, N31109, N31108, N31107, N31106, N31105, 
        N31104, N31103, N31102, N31101, N31100, N31099, N31098, N31097, N31096, 
        N31095, N31094, N31093, N31092, N31091, N31090, N31089, N31088, N31087, 
        N31086, N31085, N31084, N31083, N31082}) );
  GSIM_DW01_add_472 add_0_root_add_0_root_add_182_8 ( .A({N31145, N31144, 
        N31143, N31142, N31141, N31140, N31139, N31138, N31137, N31136, N31135, 
        N31134, N31133, N31132, N31131, N31130, N31129, N31128, N31127, N31126, 
        N31125, N31124, N31123, N31122, N31121, N31120, N31119, N31118, N31117, 
        N31116, N31115, N31114, N31113, N31112, N31111, N31110, N31109, N31108, 
        N31107, N31106, N31105, N31104, N31103, N31102, N31101, N31100, N31099, 
        N31098, N31097, N31096, N31095, N31094, N31093, N31092, N31091, N31090, 
        N31089, N31088, N31087, N31086, N31085, N31084, N31083, N31082}), .B({
        N34089, N34088, N34087, N34086, N34085, N34084, N34083, N34082, N34081, 
        N34080, N34079, N34078, N34077, N34076, N34075, N34074, N34073, N34072, 
        N34071, N34070, N34069, N34068, N34067, N34066, N34065, N34064, N34063, 
        N34062, N34061, N34060, N34059, N34058, N34057, N34056, N34055, N34054, 
        N34053, N34052, N34051, N34050, N34049, N34048, N34047, N34046, N34045, 
        N34044, N34043, N34042, N34041, N34040, N34039, N34038, N34037, N34036, 
        N34035, N34034, N34033, N34032, N34031, N34030, N34029, N34028, N34027, 
        N34026}), .CI(1'b0), .SUM({N31337, N31336, N31335, N31334, N31333, 
        N31332, N31331, N31330, N31329, N31328, N31327, N31326, N31325, N31324, 
        N31323, N31322, N31321, N31320, N31319, N31318, N31317, N31316, N31315, 
        N31314, N31313, N31312, N31311, N31310, N31309, N31308, N31307, N31306, 
        N31305, N31304, N31303, N31302, N31301, N31300, N31299, N31298, N31297, 
        N31296, N31295, N31294, N31293, N31292, N31291, N31290, N31289, N31288, 
        N31287, N31286, N31285, N31284, N31283, N31282, N31281, N31280, N31279, 
        N31278, N31277, N31276, N31275, N31274}) );
  GSIM_DW_mult_tc_8 mult_179 ( .a({1'b0, 1'b1, 1'b1, 1'b0, 1'b1}), .b({N33897, 
        N33896, N33895, N33894, N33893, N33892, N33891, N33890, N33889, N33888, 
        N33887, N33886, N33885, N33884, N33883, N33882, N33881, N33880, N33879, 
        N33878, N33877, N33876, N33875, N33874, N33873, N33872, N33871, N33870, 
        N33869, N33868, N33867, N33866, N33865, N33864, N33863, N33862, N33861, 
        N33860, N33859, N33858, N33857, N33856, N33855, N33854, N33853, N33852, 
        N33851, N33850, N33849, N33848, N33847, N33846, N33845, N33844, N33843, 
        N33842, N33841, N33840, N33839, N33838, N33837, N33836, N33835, N33834}), .product({SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, N29993, N29992, N29991, N29990, N29989, 
        N29988, N29987, N29986, N29985, N29984, N29983, N29982, N29981, N29980, 
        N29979, N29978, N29977, N29976, N29975, N29974, N29973, N29972, N29971, 
        N29970, N29969, N29968, N29967, N29966, N29965, N29964, N29963, N29962, 
        N29961, N29960, N29959, N29958, N29957, N29956, N29955, N29954, N29953, 
        N29952, N29951, N29950, N29949, N29948, N29947, N29946, N29945, N29944, 
        N29943, N29942, N29941, N29940, N29939, N29938, N29937, N29936, N29935, 
        N29934, N29933, N29932, N29931, N29930}) );
  GSIM_DW_mult_tc_7 mult_179_2 ( .a({1'b0, 1'b1, 1'b1, 1'b0, 1'b1}), .b({
        N33961, N33960, N33959, N33958, N33957, N33956, N33955, N33954, N33953, 
        N33952, N33951, N33950, N33949, N33948, N33947, N33946, N33945, N33944, 
        N33943, N33942, N33941, N33940, N33939, N33938, N33937, N33936, N33935, 
        N33934, N33933, N33932, N33931, N33930, N33929, N33928, N33927, N33926, 
        N33925, N33924, N33923, N33922, N33921, N33920, N33919, N33918, N33917, 
        N33916, N33915, N33914, N33913, N33912, N33911, N33910, N33909, N33908, 
        N33907, N33906, N33905, N33904, N33903, N33902, N33901, N33900, N33899, 
        N33898}), .product({SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, N30121, N30120, N30119, N30118, N30117, 
        N30116, N30115, N30114, N30113, N30112, N30111, N30110, N30109, N30108, 
        N30107, N30106, N30105, N30104, N30103, N30102, N30101, N30100, N30099, 
        N30098, N30097, N30096, N30095, N30094, N30093, N30092, N30091, N30090, 
        N30089, N30088, N30087, N30086, N30085, N30084, N30083, N30082, N30081, 
        N30080, N30079, N30078, N30077, N30076, N30075, N30074, N30073, N30072, 
        N30071, N30070, N30069, N30068, N30067, N30066, N30065, N30064, N30063, 
        N30062, N30061, N30060, N30059, N30058}) );
  GSIM_DW_mult_tc_6 mult_179_3 ( .a({1'b1, 1'b0, 1'b1, 1'b0}), .b({N34025, 
        N34024, N34023, N34022, N34021, N34020, N34019, N34018, N34017, N34016, 
        N34015, N34014, N34013, N34012, N34011, N34010, N34009, N34008, N34007, 
        N34006, N34005, N34004, N34003, N34002, N34001, N34000, N33999, N33998, 
        N33997, N33996, N33995, N33994, N33993, N33992, N33991, N33990, N33989, 
        N33988, N33987, N33986, N33985, N33984, N33983, N33982, N33981, N33980, 
        N33979, N33978, N33977, N33976, N33975, N33974, N33973, N33972, N33971, 
        N33970, N33969, N33968, N33967, N33966, N33965, N33964, N33963, N33962}), .product({SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, N30249, N30248, 
        N30247, N30246, N30245, N30244, N30243, N30242, N30241, N30240, N30239, 
        N30238, N30237, N30236, N30235, N30234, N30233, N30232, N30231, N30230, 
        N30229, N30228, N30227, N30226, N30225, N30224, N30223, N30222, N30221, 
        N30220, N30219, N30218, N30217, N30216, N30215, N30214, N30213, N30212, 
        N30211, N30210, N30209, N30208, N30207, N30206, N30205, N30204, N30203, 
        N30202, N30201, N30200, N30199, N30198, N30197, N30196, N30195, N30194, 
        N30193, N30192, N30191, N30190, N30189, N30188, N30187, 
        SYNOPSYS_UNCONNECTED__59}) );
  GSIM_DW01_add_483 add_3_root_add_0_root_add_179_7 ( .A({N28833, N28834, 
        N28835, N28836, N28837, N28838, N28839, N28840, N28841, N28842, N28843, 
        N28844, N28845, N28846, N28847, N28848, N28849, N28850, N28851, N28852, 
        N28853, N28854, N28855, N28856, N28857, N28858, N28859, N28860, N28861, 
        N28862, N28863, N28864, N28865, N28866, N28867, N28868, N28869, N28870, 
        N28871, N28872, N28873, N28874, N28875, N28876, N28877, N28878, N28879, 
        N28880, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N30249, N30248, N30247, 
        N30246, N30245, N30244, N30243, N30242, N30241, N30240, N30239, N30238, 
        N30237, N30236, N30235, N30234, N30233, N30232, N30231, N30230, N30229, 
        N30228, N30227, N30226, N30225, N30224, N30223, N30222, N30221, N30220, 
        N30219, N30218, N30217, N30216, N30215, N30214, N30213, N30212, N30211, 
        N30210, N30209, N30208, N30207, N30206, N30205, N30204, N30203, N30202, 
        N30201, N30200, N30199, N30198, N30197, N30196, N30195, N30194, N30193, 
        N30192, N30191, N30190, N30189, N30188, N30187, 1'b0}), .CI(1'b0), 
        .SUM({N30057, N30056, N30055, N30054, N30053, N30052, N30051, N30050, 
        N30049, N30048, N30047, N30046, N30045, N30044, N30043, N30042, N30041, 
        N30040, N30039, N30038, N30037, N30036, N30035, N30034, N30033, N30032, 
        N30031, N30030, N30029, N30028, N30027, N30026, N30025, N30024, N30023, 
        N30022, N30021, N30020, N30019, N30018, N30017, N30016, N30015, N30014, 
        N30013, N30012, N30011, N30010, N30009, N30008, N30007, N30006, N30005, 
        N30004, N30003, N30002, N30001, N30000, N29999, N29998, N29997, N29996, 
        N29995, SYNOPSYS_UNCONNECTED__60}) );
  GSIM_DW01_add_482 add_2_root_add_0_root_add_179_7 ( .A({N30057, N30056, 
        N30055, N30054, N30053, N30052, N30051, N30050, N30049, N30048, N30047, 
        N30046, N30045, N30044, N30043, N30042, N30041, N30040, N30039, N30038, 
        N30037, N30036, N30035, N30034, N30033, N30032, N30031, N30030, N30029, 
        N30028, N30027, N30026, N30025, N30024, N30023, N30022, N30021, N30020, 
        N30019, N30018, N30017, N30016, N30015, N30014, N30013, N30012, N30011, 
        N30010, N30009, N30008, N30007, N30006, N30005, N30004, N30003, N30002, 
        N30001, N30000, N29999, N29998, N29997, N29996, N29995, 1'b0}), .B({
        N29993, N29992, N29991, N29990, N29989, N29988, N29987, N29986, N29985, 
        N29984, N29983, N29982, N29981, N29980, N29979, N29978, N29977, N29976, 
        N29975, N29974, N29973, N29972, N29971, N29970, N29969, N29968, N29967, 
        N29966, N29965, N29964, N29963, N29962, N29961, N29960, N29959, N29958, 
        N29957, N29956, N29955, N29954, N29953, N29952, N29951, N29950, N29949, 
        N29948, N29947, N29946, N29945, N29944, N29943, N29942, N29941, N29940, 
        N29939, N29938, N29937, N29936, N29935, N29934, N29933, N29932, N29931, 
        N29930}), .CI(1'b0), .SUM({N30313, N30312, N30311, N30310, N30309, 
        N30308, N30307, N30306, N30305, N30304, N30303, N30302, N30301, N30300, 
        N30299, N30298, N30297, N30296, N30295, N30294, N30293, N30292, N30291, 
        N30290, N30289, N30288, N30287, N30286, N30285, N30284, N30283, N30282, 
        N30281, N30280, N30279, N30278, N30277, N30276, N30275, N30274, N30273, 
        N30272, N30271, N30270, N30269, N30268, N30267, N30266, N30265, N30264, 
        N30263, N30262, N30261, N30260, N30259, N30258, N30257, N30256, N30255, 
        N30254, N30253, N30252, N30251, N30250}) );
  GSIM_DW01_add_481 add_1_root_add_0_root_add_179_7 ( .A({N30121, N30120, 
        N30119, N30118, N30117, N30116, N30115, N30114, N30113, N30112, N30111, 
        N30110, N30109, N30108, N30107, N30106, N30105, N30104, N30103, N30102, 
        N30101, N30100, N30099, N30098, N30097, N30096, N30095, N30094, N30093, 
        N30092, N30091, N30090, N30089, N30088, N30087, N30086, N30085, N30084, 
        N30083, N30082, N30081, N30080, N30079, N30078, N30077, N30076, N30075, 
        N30074, N30073, N30072, N30071, N30070, N30069, N30068, N30067, N30066, 
        N30065, N30064, N30063, N30062, N30061, N30060, N30059, N30058}), .B({
        N30313, N30312, N30311, N30310, N30309, N30308, N30307, N30306, N30305, 
        N30304, N30303, N30302, N30301, N30300, N30299, N30298, N30297, N30296, 
        N30295, N30294, N30293, N30292, N30291, N30290, N30289, N30288, N30287, 
        N30286, N30285, N30284, N30283, N30282, N30281, N30280, N30279, N30278, 
        N30277, N30276, N30275, N30274, N30273, N30272, N30271, N30270, N30269, 
        N30268, N30267, N30266, N30265, N30264, N30263, N30262, N30261, N30260, 
        N30259, N30258, N30257, N30256, N30255, N30254, N30253, N30252, N30251, 
        N30250}), .CI(1'b0), .SUM({N30185, N30184, N30183, N30182, N30181, 
        N30180, N30179, N30178, N30177, N30176, N30175, N30174, N30173, N30172, 
        N30171, N30170, N30169, N30168, N30167, N30166, N30165, N30164, N30163, 
        N30162, N30161, N30160, N30159, N30158, N30157, N30156, N30155, N30154, 
        N30153, N30152, N30151, N30150, N30149, N30148, N30147, N30146, N30145, 
        N30144, N30143, N30142, N30141, N30140, N30139, N30138, N30137, N30136, 
        N30135, N30134, N30133, N30132, N30131, N30130, N30129, N30128, N30127, 
        N30126, N30125, N30124, N30123, N30122}) );
  GSIM_DW01_add_480 add_0_root_add_0_root_add_179_7 ( .A({N30185, N30184, 
        N30183, N30182, N30181, N30180, N30179, N30178, N30177, N30176, N30175, 
        N30174, N30173, N30172, N30171, N30170, N30169, N30168, N30167, N30166, 
        N30165, N30164, N30163, N30162, N30161, N30160, N30159, N30158, N30157, 
        N30156, N30155, N30154, N30153, N30152, N30151, N30150, N30149, N30148, 
        N30147, N30146, N30145, N30144, N30143, N30142, N30141, N30140, N30139, 
        N30138, N30137, N30136, N30135, N30134, N30133, N30132, N30131, N30130, 
        N30129, N30128, N30127, N30126, N30125, N30124, N30123, N30122}), .B({
        N34089, N34088, N34087, N34086, N34085, N34084, N34083, N34082, N34081, 
        N34080, N34079, N34078, N34077, N34076, N34075, N34074, N34073, N34072, 
        N34071, N34070, N34069, N34068, N34067, N34066, N34065, N34064, N34063, 
        N34062, N34061, N34060, N34059, N34058, N34057, N34056, N34055, N34054, 
        N34053, N34052, N34051, N34050, N34049, N34048, N34047, N34046, N34045, 
        N34044, N34043, N34042, N34041, N34040, N34039, N34038, N34037, N34036, 
        N34035, N34034, N34033, N34032, N34031, N34030, N34029, N34028, N34027, 
        N34026}), .CI(1'b0), .SUM({N30377, N30376, N30375, N30374, N30373, 
        N30372, N30371, N30370, N30369, N30368, N30367, N30366, N30365, N30364, 
        N30363, N30362, N30361, N30360, N30359, N30358, N30357, N30356, N30355, 
        N30354, N30353, N30352, N30351, N30350, N30349, N30348, N30347, N30346, 
        N30345, N30344, N30343, N30342, N30341, N30340, N30339, N30338, N30337, 
        N30336, N30335, N30334, N30333, N30332, N30331, N30330, N30329, N30328, 
        N30327, N30326, N30325, N30324, N30323, N30322, N30321, N30320, N30319, 
        N30318, N30317, N30316, N30315, N30314}) );
  GSIM_DW_mult_tc_12 mult_191_2 ( .a({1'b1, 1'b0, 1'b1, 1'b0}), .b({N33833, 
        N33832, N33831, N33830, N33829, N33828, N33827, N33826, N33825, N33824, 
        N33823, N33822, N33821, N33820, N33819, N33818, N33817, N33816, N33815, 
        N33814, N33813, N33812, N33811, N33810, N33809, N33808, N33807, N33806, 
        N33805, N33804, N33803, N33802, N33801, N33800, N33799, N33798, N33797, 
        N33796, N33795, N33794, N33793, N33792, N33791, N33790, N33789, N33788, 
        N33787, N33786, N33785, N33784, N33783, N33782, N33781, N33780, N33779, 
        N33778, N33777, N33776, N33775, N33774, N33773, N33772, N33771, N33770}), .product({SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, 
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, N33193, N33192, 
        N33191, N33190, N33189, N33188, N33187, N33186, N33185, N33184, N33183, 
        N33182, N33181, N33180, N33179, N33178, N33177, N33176, N33175, N33174, 
        N33173, N33172, N33171, N33170, N33169, N33168, N33167, N33166, N33165, 
        N33164, N33163, N33162, N33161, N33160, N33159, N33158, N33157, N33156, 
        N33155, N33154, N33153, N33152, N33151, N33150, N33149, N33148, N33147, 
        N33146, N33145, N33144, N33143, N33142, N33141, N33140, N33139, N33138, 
        N33137, N33136, N33135, N33134, N33133, N33132, N33131, 
        SYNOPSYS_UNCONNECTED__65}) );
  GSIM_DW01_add_488 add_4_root_add_0_root_add_191_7 ( .A({N28833, N28834, 
        N28835, N28836, N28837, N28838, N28839, N28840, N28841, N28842, N28843, 
        N28844, N28845, N28846, N28847, N28848, N28849, N28850, N28851, N28852, 
        N28853, N28854, N28855, N28856, N28857, N28858, N28859, N28860, N28861, 
        N28862, N28863, N28864, N28865, N28866, N28867, N28868, N28869, N28870, 
        N28871, N28872, N28873, N28874, N28875, N28876, N28877, N28878, N28879, 
        N28880, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N33193, N33192, N33191, 
        N33190, N33189, N33188, N33187, N33186, N33185, N33184, N33183, N33182, 
        N33181, N33180, N33179, N33178, N33177, N33176, N33175, N33174, N33173, 
        N33172, N33171, N33170, N33169, N33168, N33167, N33166, N33165, N33164, 
        N33163, N33162, N33161, N33160, N33159, N33158, N33157, N33156, N33155, 
        N33154, N33153, N33152, N33151, N33150, N33149, N33148, N33147, N33146, 
        N33145, N33144, N33143, N33142, N33141, N33140, N33139, N33138, N33137, 
        N33136, N33135, N33134, N33133, N33132, N33131, 1'b0}), .CI(1'b0), 
        .SUM({N33257, N33256, N33255, N33254, N33253, N33252, N33251, N33250, 
        N33249, N33248, N33247, N33246, N33245, N33244, N33243, N33242, N33241, 
        N33240, N33239, N33238, N33237, N33236, N33235, N33234, N33233, N33232, 
        N33231, N33230, N33229, N33228, N33227, N33226, N33225, N33224, N33223, 
        N33222, N33221, N33220, N33219, N33218, N33217, N33216, N33215, N33214, 
        N33213, N33212, N33211, N33210, N33209, N33208, N33207, N33206, N33205, 
        N33204, N33203, N33202, N33201, N33200, N33199, N33198, N33197, N33196, 
        N33195, SYNOPSYS_UNCONNECTED__66}) );
  GSIM_DW_mult_tc_11 mult_191_5 ( .a({1'b1, 1'b0, 1'b1, 1'b0}), .b({N34025, 
        N34024, N34023, N34022, N34021, N34020, N34019, N34018, N34017, N34016, 
        N34015, N34014, N34013, N34012, N34011, N34010, N34009, N34008, N34007, 
        N34006, N34005, N34004, N34003, N34002, N34001, N34000, N33999, N33998, 
        N33997, N33996, N33995, N33994, N33993, N33992, N33991, N33990, N33989, 
        N33988, N33987, N33986, N33985, N33984, N33983, N33982, N33981, N33980, 
        N33979, N33978, N33977, N33976, N33975, N33974, N33973, N33972, N33971, 
        N33970, N33969, N33968, N33967, N33966, N33965, N33964, N33963, N33962}), .product({SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, N33577, N33576, 
        N33575, N33574, N33573, N33572, N33571, N33570, N33569, N33568, N33567, 
        N33566, N33565, N33564, N33563, N33562, N33561, N33560, N33559, N33558, 
        N33557, N33556, N33555, N33554, N33553, N33552, N33551, N33550, N33549, 
        N33548, N33547, N33546, N33545, N33544, N33543, N33542, N33541, N33540, 
        N33539, N33538, N33537, N33536, N33535, N33534, N33533, N33532, N33531, 
        N33530, N33529, N33528, N33527, N33526, N33525, N33524, N33523, N33522, 
        N33521, N33520, N33519, N33518, N33517, N33516, N33515, 
        SYNOPSYS_UNCONNECTED__71}) );
  GSIM_DW01_add_487 add_3_root_add_0_root_add_191_7 ( .A({N33257, N33256, 
        N33255, N33254, N33253, N33252, N33251, N33250, N33249, N33248, N33247, 
        N33246, N33245, N33244, N33243, N33242, N33241, N33240, N33239, N33238, 
        N33237, N33236, N33235, N33234, N33233, N33232, N33231, N33230, N33229, 
        N33228, N33227, N33226, N33225, N33224, N33223, N33222, N33221, N33220, 
        N33219, N33218, N33217, N33216, N33215, N33214, N33213, N33212, N33211, 
        N33210, N33209, N33208, N33207, N33206, N33205, N33204, N33203, N33202, 
        N33201, N33200, N33199, N33198, N33197, N33196, N33195, 1'b0}), .B({
        N33577, N33576, N33575, N33574, N33573, N33572, N33571, N33570, N33569, 
        N33568, N33567, N33566, N33565, N33564, N33563, N33562, N33561, N33560, 
        N33559, N33558, N33557, N33556, N33555, N33554, N33553, N33552, N33551, 
        N33550, N33549, N33548, N33547, N33546, N33545, N33544, N33543, N33542, 
        N33541, N33540, N33539, N33538, N33537, N33536, N33535, N33534, N33533, 
        N33532, N33531, N33530, N33529, N33528, N33527, N33526, N33525, N33524, 
        N33523, N33522, N33521, N33520, N33519, N33518, N33517, N33516, N33515, 
        1'b0}), .CI(1'b0), .SUM({N33129, N33128, N33127, N33126, N33125, 
        N33124, N33123, N33122, N33121, N33120, N33119, N33118, N33117, N33116, 
        N33115, N33114, N33113, N33112, N33111, N33110, N33109, N33108, N33107, 
        N33106, N33105, N33104, N33103, N33102, N33101, N33100, N33099, N33098, 
        N33097, N33096, N33095, N33094, N33093, N33092, N33091, N33090, N33089, 
        N33088, N33087, N33086, N33085, N33084, N33083, N33082, N33081, N33080, 
        N33079, N33078, N33077, N33076, N33075, N33074, N33073, N33072, N33071, 
        N33070, N33069, N33068, N33067, SYNOPSYS_UNCONNECTED__72}) );
  GSIM_DW_mult_tc_10 mult_191_3 ( .a({1'b0, 1'b1, 1'b1, 1'b0, 1'b1}), .b({
        N33897, N33896, N33895, N33894, N33893, N33892, N33891, N33890, N33889, 
        N33888, N33887, N33886, N33885, N33884, N33883, N33882, N33881, N33880, 
        N33879, N33878, N33877, N33876, N33875, N33874, N33873, N33872, N33871, 
        N33870, N33869, N33868, N33867, N33866, N33865, N33864, N33863, N33862, 
        N33861, N33860, N33859, N33858, N33857, N33856, N33855, N33854, N33853, 
        N33852, N33851, N33850, N33849, N33848, N33847, N33846, N33845, N33844, 
        N33843, N33842, N33841, N33840, N33839, N33838, N33837, N33836, N33835, 
        N33834}), .product({SYNOPSYS_UNCONNECTED__73, SYNOPSYS_UNCONNECTED__74, 
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, N33321, N33320, N33319, N33318, N33317, 
        N33316, N33315, N33314, N33313, N33312, N33311, N33310, N33309, N33308, 
        N33307, N33306, N33305, N33304, N33303, N33302, N33301, N33300, N33299, 
        N33298, N33297, N33296, N33295, N33294, N33293, N33292, N33291, N33290, 
        N33289, N33288, N33287, N33286, N33285, N33284, N33283, N33282, N33281, 
        N33280, N33279, N33278, N33277, N33276, N33275, N33274, N33273, N33272, 
        N33271, N33270, N33269, N33268, N33267, N33266, N33265, N33264, N33263, 
        N33262, N33261, N33260, N33259, N33258}) );
  GSIM_DW_mult_tc_9 mult_191_4 ( .a({1'b0, 1'b1, 1'b1, 1'b0, 1'b1}), .b({
        N33961, N33960, N33959, N33958, N33957, N33956, N33955, N33954, N33953, 
        N33952, N33951, N33950, N33949, N33948, N33947, N33946, N33945, N33944, 
        N33943, N33942, N33941, N33940, N33939, N33938, N33937, N33936, N33935, 
        N33934, N33933, N33932, N33931, N33930, N33929, N33928, N33927, N33926, 
        N33925, N33924, N33923, N33922, N33921, N33920, N33919, N33918, N33917, 
        N33916, N33915, N33914, N33913, N33912, N33911, N33910, N33909, N33908, 
        N33907, N33906, N33905, N33904, N33903, N33902, N33901, N33900, N33899, 
        N33898}), .product({SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, N33449, N33448, N33447, N33446, N33445, 
        N33444, N33443, N33442, N33441, N33440, N33439, N33438, N33437, N33436, 
        N33435, N33434, N33433, N33432, N33431, N33430, N33429, N33428, N33427, 
        N33426, N33425, N33424, N33423, N33422, N33421, N33420, N33419, N33418, 
        N33417, N33416, N33415, N33414, N33413, N33412, N33411, N33410, N33409, 
        N33408, N33407, N33406, N33405, N33404, N33403, N33402, N33401, N33400, 
        N33399, N33398, N33397, N33396, N33395, N33394, N33393, N33392, N33391, 
        N33390, N33389, N33388, N33387, N33386}) );
  GSIM_DW01_add_486 add_2_root_add_0_root_add_191_7 ( .A({N33129, N33128, 
        N33127, N33126, N33125, N33124, N33123, N33122, N33121, N33120, N33119, 
        N33118, N33117, N33116, N33115, N33114, N33113, N33112, N33111, N33110, 
        N33109, N33108, N33107, N33106, N33105, N33104, N33103, N33102, N33101, 
        N33100, N33099, N33098, N33097, N33096, N33095, N33094, N33093, N33092, 
        N33091, N33090, N33089, N33088, N33087, N33086, N33085, N33084, N33083, 
        N33082, N33081, N33080, N33079, N33078, N33077, N33076, N33075, N33074, 
        N33073, N33072, N33071, N33070, N33069, N33068, N33067, 1'b0}), .B({
        N33321, N33320, N33319, N33318, N33317, N33316, N33315, N33314, N33313, 
        N33312, N33311, N33310, N33309, N33308, N33307, N33306, N33305, N33304, 
        N33303, N33302, N33301, N33300, N33299, N33298, N33297, N33296, N33295, 
        N33294, N33293, N33292, N33291, N33290, N33289, N33288, N33287, N33286, 
        N33285, N33284, N33283, N33282, N33281, N33280, N33279, N33278, N33277, 
        N33276, N33275, N33274, N33273, N33272, N33271, N33270, N33269, N33268, 
        N33267, N33266, N33265, N33264, N33263, N33262, N33261, N33260, N33259, 
        N33258}), .CI(1'b0), .SUM({N33513, N33512, N33511, N33510, N33509, 
        N33508, N33507, N33506, N33505, N33504, N33503, N33502, N33501, N33500, 
        N33499, N33498, N33497, N33496, N33495, N33494, N33493, N33492, N33491, 
        N33490, N33489, N33488, N33487, N33486, N33485, N33484, N33483, N33482, 
        N33481, N33480, N33479, N33478, N33477, N33476, N33475, N33474, N33473, 
        N33472, N33471, N33470, N33469, N33468, N33467, N33466, N33465, N33464, 
        N33463, N33462, N33461, N33460, N33459, N33458, N33457, N33456, N33455, 
        N33454, N33453, N33452, N33451, N33450}) );
  GSIM_DW01_add_485 add_1_root_add_0_root_add_191_7 ( .A({N33449, N33448, 
        N33447, N33446, N33445, N33444, N33443, N33442, N33441, N33440, N33439, 
        N33438, N33437, N33436, N33435, N33434, N33433, N33432, N33431, N33430, 
        N33429, N33428, N33427, N33426, N33425, N33424, N33423, N33422, N33421, 
        N33420, N33419, N33418, N33417, N33416, N33415, N33414, N33413, N33412, 
        N33411, N33410, N33409, N33408, N33407, N33406, N33405, N33404, N33403, 
        N33402, N33401, N33400, N33399, N33398, N33397, N33396, N33395, N33394, 
        N33393, N33392, N33391, N33390, N33389, N33388, N33387, N33386}), .B({
        N33513, N33512, N33511, N33510, N33509, N33508, N33507, N33506, N33505, 
        N33504, N33503, N33502, N33501, N33500, N33499, N33498, N33497, N33496, 
        N33495, N33494, N33493, N33492, N33491, N33490, N33489, N33488, N33487, 
        N33486, N33485, N33484, N33483, N33482, N33481, N33480, N33479, N33478, 
        N33477, N33476, N33475, N33474, N33473, N33472, N33471, N33470, N33469, 
        N33468, N33467, N33466, N33465, N33464, N33463, N33462, N33461, N33460, 
        N33459, N33458, N33457, N33456, N33455, N33454, N33453, N33452, N33451, 
        N33450}), .CI(1'b0), .SUM({N33385, N33384, N33383, N33382, N33381, 
        N33380, N33379, N33378, N33377, N33376, N33375, N33374, N33373, N33372, 
        N33371, N33370, N33369, N33368, N33367, N33366, N33365, N33364, N33363, 
        N33362, N33361, N33360, N33359, N33358, N33357, N33356, N33355, N33354, 
        N33353, N33352, N33351, N33350, N33349, N33348, N33347, N33346, N33345, 
        N33344, N33343, N33342, N33341, N33340, N33339, N33338, N33337, N33336, 
        N33335, N33334, N33333, N33332, N33331, N33330, N33329, N33328, N33327, 
        N33326, N33325, N33324, N33323, N33322}) );
  GSIM_DW01_add_484 add_0_root_add_0_root_add_191_7 ( .A({N33385, N33384, 
        N33383, N33382, N33381, N33380, N33379, N33378, N33377, N33376, N33375, 
        N33374, N33373, N33372, N33371, N33370, N33369, N33368, N33367, N33366, 
        N33365, N33364, N33363, N33362, N33361, N33360, N33359, N33358, N33357, 
        N33356, N33355, N33354, N33353, N33352, N33351, N33350, N33349, N33348, 
        N33347, N33346, N33345, N33344, N33343, N33342, N33341, N33340, N33339, 
        N33338, N33337, N33336, N33335, N33334, N33333, N33332, N33331, N33330, 
        N33329, N33328, N33327, N33326, N33325, N33324, N33323, N33322}), .B({
        N33769, N33768, N33767, N33766, N33765, N33764, N33763, N33762, N33761, 
        N33760, N33759, N33758, N33757, N33756, N33755, N33754, N33753, N33752, 
        N33751, N33750, N33749, N33748, N33747, N33746, N33745, N33744, N33743, 
        N33742, N33741, N33740, N33739, N33738, N33737, N33736, N33735, N33734, 
        N33733, N33732, N33731, N33730, N33729, N33728, N33727, N33726, N33725, 
        N33724, N33723, N33722, N33721, N33720, N33719, N33718, N33717, N33716, 
        N33715, N33714, N33713, N33712, N33711, N33710, N33709, N33708, N33707, 
        N33706}), .CI(1'b0), .SUM({N33641, N33640, N33639, N33638, N33637, 
        N33636, N33635, N33634, N33633, N33632, N33631, N33630, N33629, N33628, 
        N33627, N33626, N33625, N33624, N33623, N33622, N33621, N33620, N33619, 
        N33618, N33617, N33616, N33615, N33614, N33613, N33612, N33611, N33610, 
        N33609, N33608, N33607, N33606, N33605, N33604, N33603, N33602, N33601, 
        N33600, N33599, N33598, N33597, N33596, N33595, N33594, N33593, N33592, 
        N33591, N33590, N33589, N33588, N33587, N33586, N33585, N33584, N33583, 
        N33582, N33581, N33580, N33579, N33578}) );
  GSIM_DW_mult_tc_17 mult_188_2 ( .a({1'b1, 1'b0, 1'b1, 1'b0}), .b({N33833, 
        N33832, N33831, N33830, N33829, N33828, N33827, N33826, N33825, N33824, 
        N33823, N33822, N33821, N33820, N33819, N33818, N33817, N33816, N33815, 
        N33814, N33813, N33812, N33811, N33810, N33809, N33808, N33807, N33806, 
        N33805, N33804, N33803, N33802, N33801, N33800, N33799, N33798, N33797, 
        N33796, N33795, N33794, N33793, N33792, N33791, N33790, N33789, N33788, 
        N33787, N33786, N33785, N33784, N33783, N33782, N33781, N33780, N33779, 
        N33778, N33777, N33776, N33775, N33774, N33773, N33772, N33771, N33770}), .product({SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, N32361, N32360, 
        N32359, N32358, N32357, N32356, N32355, N32354, N32353, N32352, N32351, 
        N32350, N32349, N32348, N32347, N32346, N32345, N32344, N32343, N32342, 
        N32341, N32340, N32339, N32338, N32337, N32336, N32335, N32334, N32333, 
        N32332, N32331, N32330, N32329, N32328, N32327, N32326, N32325, N32324, 
        N32323, N32322, N32321, N32320, N32319, N32318, N32317, N32316, N32315, 
        N32314, N32313, N32312, N32311, N32310, N32309, N32308, N32307, N32306, 
        N32305, N32304, N32303, N32302, N32301, N32300, N32299, 
        SYNOPSYS_UNCONNECTED__87}) );
  GSIM_DW01_add_495 add_3_root_add_0_root_add_188_5 ( .A({N28833, N28834, 
        N28835, N28836, N28837, N28838, N28839, N28840, N28841, N28842, N28843, 
        N28844, N28845, N28846, N28847, N28848, N28849, N28850, N28851, N28852, 
        N28853, N28854, N28855, N28856, N28857, N28858, N28859, N28860, N28861, 
        N28862, N28863, N28864, N28865, N28866, N28867, N28868, N28869, N28870, 
        N28871, N28872, N28873, N28874, N28875, N28876, N28877, N28878, N28879, 
        N28880, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N32361, N32360, N32359, 
        N32358, N32357, N32356, N32355, N32354, N32353, N32352, N32351, N32350, 
        N32349, N32348, N32347, N32346, N32345, N32344, N32343, N32342, N32341, 
        N32340, N32339, N32338, N32337, N32336, N32335, N32334, N32333, N32332, 
        N32331, N32330, N32329, N32328, N32327, N32326, N32325, N32324, N32323, 
        N32322, N32321, N32320, N32319, N32318, N32317, N32316, N32315, N32314, 
        N32313, N32312, N32311, N32310, N32309, N32308, N32307, N32306, N32305, 
        N32304, N32303, N32302, N32301, N32300, N32299, 1'b0}), .CI(1'b0), 
        .SUM({N32297, N32296, N32295, N32294, N32293, N32292, N32291, N32290, 
        N32289, N32288, N32287, N32286, N32285, N32284, N32283, N32282, N32281, 
        N32280, N32279, N32278, N32277, N32276, N32275, N32274, N32273, N32272, 
        N32271, N32270, N32269, N32268, N32267, N32266, N32265, N32264, N32263, 
        N32262, N32261, N32260, N32259, N32258, N32257, N32256, N32255, N32254, 
        N32253, N32252, N32251, N32250, N32249, N32248, N32247, N32246, N32245, 
        N32244, N32243, N32242, N32241, N32240, N32239, N32238, N32237, N32236, 
        N32235, SYNOPSYS_UNCONNECTED__88}) );
  GSIM_DW_mult_tc_16 mult_188_3 ( .a({1'b0, 1'b1, 1'b1, 1'b0, 1'b1}), .b({
        N33897, N33896, N33895, N33894, N33893, N33892, N33891, N33890, N33889, 
        N33888, N33887, N33886, N33885, N33884, N33883, N33882, N33881, N33880, 
        N33879, N33878, N33877, N33876, N33875, N33874, N33873, N33872, N33871, 
        N33870, N33869, N33868, N33867, N33866, N33865, N33864, N33863, N33862, 
        N33861, N33860, N33859, N33858, N33857, N33856, N33855, N33854, N33853, 
        N33852, N33851, N33850, N33849, N33848, N33847, N33846, N33845, N33844, 
        N33843, N33842, N33841, N33840, N33839, N33838, N33837, N33836, N33835, 
        N33834}), .product({SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, 
        SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, 
        SYNOPSYS_UNCONNECTED__93, N32489, N32488, N32487, N32486, N32485, 
        N32484, N32483, N32482, N32481, N32480, N32479, N32478, N32477, N32476, 
        N32475, N32474, N32473, N32472, N32471, N32470, N32469, N32468, N32467, 
        N32466, N32465, N32464, N32463, N32462, N32461, N32460, N32459, N32458, 
        N32457, N32456, N32455, N32454, N32453, N32452, N32451, N32450, N32449, 
        N32448, N32447, N32446, N32445, N32444, N32443, N32442, N32441, N32440, 
        N32439, N32438, N32437, N32436, N32435, N32434, N32433, N32432, N32431, 
        N32430, N32429, N32428, N32427, N32426}) );
  GSIM_DW_mult_tc_15 mult_188_4 ( .a({1'b0, 1'b1, 1'b1, 1'b0, 1'b1}), .b({
        N33961, N33960, N33959, N33958, N33957, N33956, N33955, N33954, N33953, 
        N33952, N33951, N33950, N33949, N33948, N33947, N33946, N33945, N33944, 
        N33943, N33942, N33941, N33940, N33939, N33938, N33937, N33936, N33935, 
        N33934, N33933, N33932, N33931, N33930, N33929, N33928, N33927, N33926, 
        N33925, N33924, N33923, N33922, N33921, N33920, N33919, N33918, N33917, 
        N33916, N33915, N33914, N33913, N33912, N33911, N33910, N33909, N33908, 
        N33907, N33906, N33905, N33904, N33903, N33902, N33901, N33900, N33899, 
        N33898}), .product({SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, N32617, N32616, N32615, N32614, N32613, 
        N32612, N32611, N32610, N32609, N32608, N32607, N32606, N32605, N32604, 
        N32603, N32602, N32601, N32600, N32599, N32598, N32597, N32596, N32595, 
        N32594, N32593, N32592, N32591, N32590, N32589, N32588, N32587, N32586, 
        N32585, N32584, N32583, N32582, N32581, N32580, N32579, N32578, N32577, 
        N32576, N32575, N32574, N32573, N32572, N32571, N32570, N32569, N32568, 
        N32567, N32566, N32565, N32564, N32563, N32562, N32561, N32560, N32559, 
        N32558, N32557, N32556, N32555, N32554}) );
  GSIM_DW01_add_494 add_2_root_add_0_root_add_188_5 ( .A({N32297, N32296, 
        N32295, N32294, N32293, N32292, N32291, N32290, N32289, N32288, N32287, 
        N32286, N32285, N32284, N32283, N32282, N32281, N32280, N32279, N32278, 
        N32277, N32276, N32275, N32274, N32273, N32272, N32271, N32270, N32269, 
        N32268, N32267, N32266, N32265, N32264, N32263, N32262, N32261, N32260, 
        N32259, N32258, N32257, N32256, N32255, N32254, N32253, N32252, N32251, 
        N32250, N32249, N32248, N32247, N32246, N32245, N32244, N32243, N32242, 
        N32241, N32240, N32239, N32238, N32237, N32236, N32235, 1'b0}), .B({
        N32617, N32616, N32615, N32614, N32613, N32612, N32611, N32610, N32609, 
        N32608, N32607, N32606, N32605, N32604, N32603, N32602, N32601, N32600, 
        N32599, N32598, N32597, N32596, N32595, N32594, N32593, N32592, N32591, 
        N32590, N32589, N32588, N32587, N32586, N32585, N32584, N32583, N32582, 
        N32581, N32580, N32579, N32578, N32577, N32576, N32575, N32574, N32573, 
        N32572, N32571, N32570, N32569, N32568, N32567, N32566, N32565, N32564, 
        N32563, N32562, N32561, N32560, N32559, N32558, N32557, N32556, N32555, 
        N32554}), .CI(1'b0), .SUM({N32553, N32552, N32551, N32550, N32549, 
        N32548, N32547, N32546, N32545, N32544, N32543, N32542, N32541, N32540, 
        N32539, N32538, N32537, N32536, N32535, N32534, N32533, N32532, N32531, 
        N32530, N32529, N32528, N32527, N32526, N32525, N32524, N32523, N32522, 
        N32521, N32520, N32519, N32518, N32517, N32516, N32515, N32514, N32513, 
        N32512, N32511, N32510, N32509, N32508, N32507, N32506, N32505, N32504, 
        N32503, N32502, N32501, N32500, N32499, N32498, N32497, N32496, N32495, 
        N32494, N32493, N32492, N32491, N32490}) );
  GSIM_DW01_add_493 add_1_root_add_0_root_add_188_5 ( .A({N32489, N32488, 
        N32487, N32486, N32485, N32484, N32483, N32482, N32481, N32480, N32479, 
        N32478, N32477, N32476, N32475, N32474, N32473, N32472, N32471, N32470, 
        N32469, N32468, N32467, N32466, N32465, N32464, N32463, N32462, N32461, 
        N32460, N32459, N32458, N32457, N32456, N32455, N32454, N32453, N32452, 
        N32451, N32450, N32449, N32448, N32447, N32446, N32445, N32444, N32443, 
        N32442, N32441, N32440, N32439, N32438, N32437, N32436, N32435, N32434, 
        N32433, N32432, N32431, N32430, N32429, N32428, N32427, N32426}), .B({
        N32553, N32552, N32551, N32550, N32549, N32548, N32547, N32546, N32545, 
        N32544, N32543, N32542, N32541, N32540, N32539, N32538, N32537, N32536, 
        N32535, N32534, N32533, N32532, N32531, N32530, N32529, N32528, N32527, 
        N32526, N32525, N32524, N32523, N32522, N32521, N32520, N32519, N32518, 
        N32517, N32516, N32515, N32514, N32513, N32512, N32511, N32510, N32509, 
        N32508, N32507, N32506, N32505, N32504, N32503, N32502, N32501, N32500, 
        N32499, N32498, N32497, N32496, N32495, N32494, N32493, N32492, N32491, 
        N32490}), .CI(1'b0), .SUM({N32425, N32424, N32423, N32422, N32421, 
        N32420, N32419, N32418, N32417, N32416, N32415, N32414, N32413, N32412, 
        N32411, N32410, N32409, N32408, N32407, N32406, N32405, N32404, N32403, 
        N32402, N32401, N32400, N32399, N32398, N32397, N32396, N32395, N32394, 
        N32393, N32392, N32391, N32390, N32389, N32388, N32387, N32386, N32385, 
        N32384, N32383, N32382, N32381, N32380, N32379, N32378, N32377, N32376, 
        N32375, N32374, N32373, N32372, N32371, N32370, N32369, N32368, N32367, 
        N32366, N32365, N32364, N32363, N32362}) );
  GSIM_DW01_add_492 add_0_root_add_0_root_add_188_5 ( .A({N32425, N32424, 
        N32423, N32422, N32421, N32420, N32419, N32418, N32417, N32416, N32415, 
        N32414, N32413, N32412, N32411, N32410, N32409, N32408, N32407, N32406, 
        N32405, N32404, N32403, N32402, N32401, N32400, N32399, N32398, N32397, 
        N32396, N32395, N32394, N32393, N32392, N32391, N32390, N32389, N32388, 
        N32387, N32386, N32385, N32384, N32383, N32382, N32381, N32380, N32379, 
        N32378, N32377, N32376, N32375, N32374, N32373, N32372, N32371, N32370, 
        N32369, N32368, N32367, N32366, N32365, N32364, N32363, N32362}), .B({
        N33769, N33768, N33767, N33766, N33765, N33764, N33763, N33762, N33761, 
        N33760, N33759, N33758, N33757, N33756, N33755, N33754, N33753, N33752, 
        N33751, N33750, N33749, N33748, N33747, N33746, N33745, N33744, N33743, 
        N33742, N33741, N33740, N33739, N33738, N33737, N33736, N33735, N33734, 
        N33733, N33732, N33731, N33730, N33729, N33728, N33727, N33726, N33725, 
        N33724, N33723, N33722, N33721, N33720, N33719, N33718, N33717, N33716, 
        N33715, N33714, N33713, N33712, N33711, N33710, N33709, N33708, N33707, 
        N33706}), .CI(1'b0), .SUM({N32681, N32680, N32679, N32678, N32677, 
        N32676, N32675, N32674, N32673, N32672, N32671, N32670, N32669, N32668, 
        N32667, N32666, N32665, N32664, N32663, N32662, N32661, N32660, N32659, 
        N32658, N32657, N32656, N32655, N32654, N32653, N32652, N32651, N32650, 
        N32649, N32648, N32647, N32646, N32645, N32644, N32643, N32642, N32641, 
        N32640, N32639, N32638, N32637, N32636, N32635, N32634, N32633, N32632, 
        N32631, N32630, N32629, N32628, N32627, N32626, N32625, N32624, N32623, 
        N32622, N32621, N32620, N32619, N32618}) );
  GSIM_DW_mult_tc_14 mult_185_2 ( .a({1'b1, 1'b0, 1'b1, 1'b0}), .b({N33833, 
        N33832, N33831, N33830, N33829, N33828, N33827, N33826, N33825, N33824, 
        N33823, N33822, N33821, N33820, N33819, N33818, N33817, N33816, N33815, 
        N33814, N33813, N33812, N33811, N33810, N33809, N33808, N33807, N33806, 
        N33805, N33804, N33803, N33802, N33801, N33800, N33799, N33798, N33797, 
        N33796, N33795, N33794, N33793, N33792, N33791, N33790, N33789, N33788, 
        N33787, N33786, N33785, N33784, N33783, N33782, N33781, N33780, N33779, 
        N33778, N33777, N33776, N33775, N33774, N33773, N33772, N33771, N33770}), .product({SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, N31721, N31720, 
        N31719, N31718, N31717, N31716, N31715, N31714, N31713, N31712, N31711, 
        N31710, N31709, N31708, N31707, N31706, N31705, N31704, N31703, N31702, 
        N31701, N31700, N31699, N31698, N31697, N31696, N31695, N31694, N31693, 
        N31692, N31691, N31690, N31689, N31688, N31687, N31686, N31685, N31684, 
        N31683, N31682, N31681, N31680, N31679, N31678, N31677, N31676, N31675, 
        N31674, N31673, N31672, N31671, N31670, N31669, N31668, N31667, N31666, 
        N31665, N31664, N31663, N31662, N31661, N31660, N31659, 
        SYNOPSYS_UNCONNECTED__103}) );
  GSIM_DW01_add_491 add_2_root_add_0_root_add_185_3 ( .A({N28833, N28834, 
        N28835, N28836, N28837, N28838, N28839, N28840, N28841, N28842, N28843, 
        N28844, N28845, N28846, N28847, N28848, N28849, N28850, N28851, N28852, 
        N28853, N28854, N28855, N28856, N28857, N28858, N28859, N28860, N28861, 
        N28862, N28863, N28864, N28865, N28866, N28867, N28868, N28869, N28870, 
        N28871, N28872, N28873, N28874, N28875, N28876, N28877, N28878, N28879, 
        N28880, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N31721, N31720, N31719, 
        N31718, N31717, N31716, N31715, N31714, N31713, N31712, N31711, N31710, 
        N31709, N31708, N31707, N31706, N31705, N31704, N31703, N31702, N31701, 
        N31700, N31699, N31698, N31697, N31696, N31695, N31694, N31693, N31692, 
        N31691, N31690, N31689, N31688, N31687, N31686, N31685, N31684, N31683, 
        N31682, N31681, N31680, N31679, N31678, N31677, N31676, N31675, N31674, 
        N31673, N31672, N31671, N31670, N31669, N31668, N31667, N31666, N31665, 
        N31664, N31663, N31662, N31661, N31660, N31659, 1'b0}), .CI(1'b0), 
        .SUM({N31785, N31784, N31783, N31782, N31781, N31780, N31779, N31778, 
        N31777, N31776, N31775, N31774, N31773, N31772, N31771, N31770, N31769, 
        N31768, N31767, N31766, N31765, N31764, N31763, N31762, N31761, N31760, 
        N31759, N31758, N31757, N31756, N31755, N31754, N31753, N31752, N31751, 
        N31750, N31749, N31748, N31747, N31746, N31745, N31744, N31743, N31742, 
        N31741, N31740, N31739, N31738, N31737, N31736, N31735, N31734, N31733, 
        N31732, N31731, N31730, N31729, N31728, N31727, N31726, N31725, N31724, 
        N31723, SYNOPSYS_UNCONNECTED__104}) );
  GSIM_DW_mult_tc_13 mult_185_3 ( .a({1'b0, 1'b1, 1'b1, 1'b0, 1'b1}), .b({
        N33897, N33896, N33895, N33894, N33893, N33892, N33891, N33890, N33889, 
        N33888, N33887, N33886, N33885, N33884, N33883, N33882, N33881, N33880, 
        N33879, N33878, N33877, N33876, N33875, N33874, N33873, N33872, N33871, 
        N33870, N33869, N33868, N33867, N33866, N33865, N33864, N33863, N33862, 
        N33861, N33860, N33859, N33858, N33857, N33856, N33855, N33854, N33853, 
        N33852, N33851, N33850, N33849, N33848, N33847, N33846, N33845, N33844, 
        N33843, N33842, N33841, N33840, N33839, N33838, N33837, N33836, N33835, 
        N33834}), .product({SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, N31849, N31848, 
        N31847, N31846, N31845, N31844, N31843, N31842, N31841, N31840, N31839, 
        N31838, N31837, N31836, N31835, N31834, N31833, N31832, N31831, N31830, 
        N31829, N31828, N31827, N31826, N31825, N31824, N31823, N31822, N31821, 
        N31820, N31819, N31818, N31817, N31816, N31815, N31814, N31813, N31812, 
        N31811, N31810, N31809, N31808, N31807, N31806, N31805, N31804, N31803, 
        N31802, N31801, N31800, N31799, N31798, N31797, N31796, N31795, N31794, 
        N31793, N31792, N31791, N31790, N31789, N31788, N31787, N31786}) );
  GSIM_DW01_add_490 add_1_root_add_0_root_add_185_3 ( .A({N31785, N31784, 
        N31783, N31782, N31781, N31780, N31779, N31778, N31777, N31776, N31775, 
        N31774, N31773, N31772, N31771, N31770, N31769, N31768, N31767, N31766, 
        N31765, N31764, N31763, N31762, N31761, N31760, N31759, N31758, N31757, 
        N31756, N31755, N31754, N31753, N31752, N31751, N31750, N31749, N31748, 
        N31747, N31746, N31745, N31744, N31743, N31742, N31741, N31740, N31739, 
        N31738, N31737, N31736, N31735, N31734, N31733, N31732, N31731, N31730, 
        N31729, N31728, N31727, N31726, N31725, N31724, N31723, 1'b0}), .B({
        N31849, N31848, N31847, N31846, N31845, N31844, N31843, N31842, N31841, 
        N31840, N31839, N31838, N31837, N31836, N31835, N31834, N31833, N31832, 
        N31831, N31830, N31829, N31828, N31827, N31826, N31825, N31824, N31823, 
        N31822, N31821, N31820, N31819, N31818, N31817, N31816, N31815, N31814, 
        N31813, N31812, N31811, N31810, N31809, N31808, N31807, N31806, N31805, 
        N31804, N31803, N31802, N31801, N31800, N31799, N31798, N31797, N31796, 
        N31795, N31794, N31793, N31792, N31791, N31790, N31789, N31788, N31787, 
        N31786}), .CI(1'b0), .SUM({N31657, N31656, N31655, N31654, N31653, 
        N31652, N31651, N31650, N31649, N31648, N31647, N31646, N31645, N31644, 
        N31643, N31642, N31641, N31640, N31639, N31638, N31637, N31636, N31635, 
        N31634, N31633, N31632, N31631, N31630, N31629, N31628, N31627, N31626, 
        N31625, N31624, N31623, N31622, N31621, N31620, N31619, N31618, N31617, 
        N31616, N31615, N31614, N31613, N31612, N31611, N31610, N31609, N31608, 
        N31607, N31606, N31605, N31604, N31603, N31602, N31601, N31600, N31599, 
        N31598, N31597, N31596, N31595, N31594}) );
  GSIM_DW01_add_489 add_0_root_add_0_root_add_185_3 ( .A({N31657, N31656, 
        N31655, N31654, N31653, N31652, N31651, N31650, N31649, N31648, N31647, 
        N31646, N31645, N31644, N31643, N31642, N31641, N31640, N31639, N31638, 
        N31637, N31636, N31635, N31634, N31633, N31632, N31631, N31630, N31629, 
        N31628, N31627, N31626, N31625, N31624, N31623, N31622, N31621, N31620, 
        N31619, N31618, N31617, N31616, N31615, N31614, N31613, N31612, N31611, 
        N31610, N31609, N31608, N31607, N31606, N31605, N31604, N31603, N31602, 
        N31601, N31600, N31599, N31598, N31597, N31596, N31595, N31594}), .B({
        N33769, N33768, N33767, N33766, N33765, N33764, N33763, N33762, N33761, 
        N33760, N33759, N33758, N33757, N33756, N33755, N33754, N33753, N33752, 
        N33751, N33750, N33749, N33748, N33747, N33746, N33745, N33744, N33743, 
        N33742, N33741, N33740, N33739, N33738, N33737, N33736, N33735, N33734, 
        N33733, N33732, N33731, N33730, N33729, N33728, N33727, N33726, N33725, 
        N33724, N33723, N33722, N33721, N33720, N33719, N33718, N33717, N33716, 
        N33715, N33714, N33713, N33712, N33711, N33710, N33709, N33708, N33707, 
        N33706}), .CI(1'b0), .SUM({N31913, N31912, N31911, N31910, N31909, 
        N31908, N31907, N31906, N31905, N31904, N31903, N31902, N31901, N31900, 
        N31899, N31898, N31897, N31896, N31895, N31894, N31893, N31892, N31891, 
        N31890, N31889, N31888, N31887, N31886, N31885, N31884, N31883, N31882, 
        N31881, N31880, N31879, N31878, N31877, N31876, N31875, N31874, N31873, 
        N31872, N31871, N31870, N31869, N31868, N31867, N31866, N31865, N31864, 
        N31863, N31862, N31861, N31860, N31859, N31858, N31857, N31856, N31855, 
        N31854, N31853, N31852, N31851, N31850}) );
  GSIM_DW_mult_tc_5 mult_176 ( .a({1'b0, 1'b1, 1'b1, 1'b0, 1'b1}), .b({N33961, 
        N33960, N33959, N33958, N33957, N33956, N33955, N33954, N33953, N33952, 
        N33951, N33950, N33949, N33948, N33947, N33946, N33945, N33944, N33943, 
        N33942, N33941, N33940, N33939, N33938, N33937, N33936, N33935, N33934, 
        N33933, N33932, N33931, N33930, N33929, N33928, N33927, N33926, N33925, 
        N33924, N33923, N33922, N33921, N33920, N33919, N33918, N33917, N33916, 
        N33915, N33914, N33913, N33912, N33911, N33910, N33909, N33908, N33907, 
        N33906, N33905, N33904, N33903, N33902, N33901, N33900, N33899, N33898}), .product({SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, N29353, N29352, N29351, N29350, N29349, 
        N29348, N29347, N29346, N29345, N29344, N29343, N29342, N29341, N29340, 
        N29339, N29338, N29337, N29336, N29335, N29334, N29333, N29332, N29331, 
        N29330, N29329, N29328, N29327, N29326, N29325, N29324, N29323, N29322, 
        N29321, N29320, N29319, N29318, N29317, N29316, N29315, N29314, N29313, 
        N29312, N29311, N29310, N29309, N29308, N29307, N29306, N29305, N29304, 
        N29303, N29302, N29301, N29300, N29299, N29298, N29297, N29296, N29295, 
        N29294, N29293, N29292, N29291, N29290}) );
  GSIM_DW_mult_tc_4 mult_176_2 ( .a({1'b1, 1'b0, 1'b1, 1'b0}), .b({N34025, 
        N34024, N34023, N34022, N34021, N34020, N34019, N34018, N34017, N34016, 
        N34015, N34014, N34013, N34012, N34011, N34010, N34009, N34008, N34007, 
        N34006, N34005, N34004, N34003, N34002, N34001, N34000, N33999, N33998, 
        N33997, N33996, N33995, N33994, N33993, N33992, N33991, N33990, N33989, 
        N33988, N33987, N33986, N33985, N33984, N33983, N33982, N33981, N33980, 
        N33979, N33978, N33977, N33976, N33975, N33974, N33973, N33972, N33971, 
        N33970, N33969, N33968, N33967, N33966, N33965, N33964, N33963, N33962}), .product({SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, N29481, N29480, 
        N29479, N29478, N29477, N29476, N29475, N29474, N29473, N29472, N29471, 
        N29470, N29469, N29468, N29467, N29466, N29465, N29464, N29463, N29462, 
        N29461, N29460, N29459, N29458, N29457, N29456, N29455, N29454, N29453, 
        N29452, N29451, N29450, N29449, N29448, N29447, N29446, N29445, N29444, 
        N29443, N29442, N29441, N29440, N29439, N29438, N29437, N29436, N29435, 
        N29434, N29433, N29432, N29431, N29430, N29429, N29428, N29427, N29426, 
        N29425, N29424, N29423, N29422, N29421, N29420, N29419, 
        SYNOPSYS_UNCONNECTED__119}) );
  GSIM_DW01_add_479 add_2_root_add_0_root_add_176_6 ( .A({N28833, N28834, 
        N28835, N28836, N28837, N28838, N28839, N28840, N28841, N28842, N28843, 
        N28844, N28845, N28846, N28847, N28848, N28849, N28850, N28851, N28852, 
        N28853, N28854, N28855, N28856, N28857, N28858, N28859, N28860, N28861, 
        N28862, N28863, N28864, N28865, N28866, N28867, N28868, N28869, N28870, 
        N28871, N28872, N28873, N28874, N28875, N28876, N28877, N28878, N28879, 
        N28880, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N29481, N29480, N29479, 
        N29478, N29477, N29476, N29475, N29474, N29473, N29472, N29471, N29470, 
        N29469, N29468, N29467, N29466, N29465, N29464, N29463, N29462, N29461, 
        N29460, N29459, N29458, N29457, N29456, N29455, N29454, N29453, N29452, 
        N29451, N29450, N29449, N29448, N29447, N29446, N29445, N29444, N29443, 
        N29442, N29441, N29440, N29439, N29438, N29437, N29436, N29435, N29434, 
        N29433, N29432, N29431, N29430, N29429, N29428, N29427, N29426, N29425, 
        N29424, N29423, N29422, N29421, N29420, N29419, 1'b0}), .CI(1'b0), 
        .SUM({N29545, N29544, N29543, N29542, N29541, N29540, N29539, N29538, 
        N29537, N29536, N29535, N29534, N29533, N29532, N29531, N29530, N29529, 
        N29528, N29527, N29526, N29525, N29524, N29523, N29522, N29521, N29520, 
        N29519, N29518, N29517, N29516, N29515, N29514, N29513, N29512, N29511, 
        N29510, N29509, N29508, N29507, N29506, N29505, N29504, N29503, N29502, 
        N29501, N29500, N29499, N29498, N29497, N29496, N29495, N29494, N29493, 
        N29492, N29491, N29490, N29489, N29488, N29487, N29486, N29485, N29484, 
        N29483, SYNOPSYS_UNCONNECTED__120}) );
  GSIM_DW01_add_478 add_1_root_add_0_root_add_176_6 ( .A({N29545, N29544, 
        N29543, N29542, N29541, N29540, N29539, N29538, N29537, N29536, N29535, 
        N29534, N29533, N29532, N29531, N29530, N29529, N29528, N29527, N29526, 
        N29525, N29524, N29523, N29522, N29521, N29520, N29519, N29518, N29517, 
        N29516, N29515, N29514, N29513, N29512, N29511, N29510, N29509, N29508, 
        N29507, N29506, N29505, N29504, N29503, N29502, N29501, N29500, N29499, 
        N29498, N29497, N29496, N29495, N29494, N29493, N29492, N29491, N29490, 
        N29489, N29488, N29487, N29486, N29485, N29484, N29483, 1'b0}), .B({
        N29353, N29352, N29351, N29350, N29349, N29348, N29347, N29346, N29345, 
        N29344, N29343, N29342, N29341, N29340, N29339, N29338, N29337, N29336, 
        N29335, N29334, N29333, N29332, N29331, N29330, N29329, N29328, N29327, 
        N29326, N29325, N29324, N29323, N29322, N29321, N29320, N29319, N29318, 
        N29317, N29316, N29315, N29314, N29313, N29312, N29311, N29310, N29309, 
        N29308, N29307, N29306, N29305, N29304, N29303, N29302, N29301, N29300, 
        N29299, N29298, N29297, N29296, N29295, N29294, N29293, N29292, N29291, 
        N29290}), .CI(1'b0), .SUM({N29417, N29416, N29415, N29414, N29413, 
        N29412, N29411, N29410, N29409, N29408, N29407, N29406, N29405, N29404, 
        N29403, N29402, N29401, N29400, N29399, N29398, N29397, N29396, N29395, 
        N29394, N29393, N29392, N29391, N29390, N29389, N29388, N29387, N29386, 
        N29385, N29384, N29383, N29382, N29381, N29380, N29379, N29378, N29377, 
        N29376, N29375, N29374, N29373, N29372, N29371, N29370, N29369, N29368, 
        N29367, N29366, N29365, N29364, N29363, N29362, N29361, N29360, N29359, 
        N29358, N29357, N29356, N29355, N29354}) );
  GSIM_DW01_add_477 add_0_root_add_0_root_add_176_6 ( .A({N29417, N29416, 
        N29415, N29414, N29413, N29412, N29411, N29410, N29409, N29408, N29407, 
        N29406, N29405, N29404, N29403, N29402, N29401, N29400, N29399, N29398, 
        N29397, N29396, N29395, N29394, N29393, N29392, N29391, N29390, N29389, 
        N29388, N29387, N29386, N29385, N29384, N29383, N29382, N29381, N29380, 
        N29379, N29378, N29377, N29376, N29375, N29374, N29373, N29372, N29371, 
        N29370, N29369, N29368, N29367, N29366, N29365, N29364, N29363, N29362, 
        N29361, N29360, N29359, N29358, N29357, N29356, N29355, N29354}), .B({
        N34089, N34088, N34087, N34086, N34085, N34084, N34083, N34082, N34081, 
        N34080, N34079, N34078, N34077, N34076, N34075, N34074, N34073, N34072, 
        N34071, N34070, N34069, N34068, N34067, N34066, N34065, N34064, N34063, 
        N34062, N34061, N34060, N34059, N34058, N34057, N34056, N34055, N34054, 
        N34053, N34052, N34051, N34050, N34049, N34048, N34047, N34046, N34045, 
        N34044, N34043, N34042, N34041, N34040, N34039, N34038, N34037, N34036, 
        N34035, N34034, N34033, N34032, N34031, N34030, N34029, N34028, N34027, 
        N34026}), .CI(1'b0), .SUM({N29609, N29608, N29607, N29606, N29605, 
        N29604, N29603, N29602, N29601, N29600, N29599, N29598, N29597, N29596, 
        N29595, N29594, N29593, N29592, N29591, N29590, N29589, N29588, N29587, 
        N29586, N29585, N29584, N29583, N29582, N29581, N29580, N29579, N29578, 
        N29577, N29576, N29575, N29574, N29573, N29572, N29571, N29570, N29569, 
        N29568, N29567, N29566, N29565, N29564, N29563, N29562, N29561, N29560, 
        N29559, N29558, N29557, N29556, N29555, N29554, N29553, N29552, N29551, 
        N29550, N29549, N29548, N29547, N29546}) );
  DFFRX1 \outCount_reg[31]  ( .D(outCount_next[31]), .CK(clk), .RN(n7647), .Q(
        outCount[31]) );
  DFFRX1 \inCount_reg[13]  ( .D(N1819), .CK(clk), .RN(n7637), .Q(inCount[13]), 
        .QN(n83) );
  DFFRX1 \inCount_reg[14]  ( .D(N1820), .CK(clk), .RN(n7637), .Q(inCount[14]), 
        .QN(n84) );
  DFFRX1 \inCount_reg[15]  ( .D(N1821), .CK(clk), .RN(n7637), .Q(inCount[15]), 
        .QN(n85) );
  DFFRX1 \inCount_reg[16]  ( .D(N1822), .CK(clk), .RN(n7638), .Q(inCount[16]), 
        .QN(n86) );
  DFFRX1 \inCount_reg[17]  ( .D(N1823), .CK(clk), .RN(n7638), .Q(inCount[17]), 
        .QN(n87) );
  DFFRX1 \inCount_reg[18]  ( .D(N1824), .CK(clk), .RN(n7638), .Q(inCount[18]), 
        .QN(n88) );
  DFFRX1 \inCount_reg[21]  ( .D(N1827), .CK(clk), .RN(n7638), .Q(inCount[21]), 
        .QN(n91) );
  DFFRX1 \inCount_reg[26]  ( .D(N1832), .CK(clk), .RN(n7638), .Q(inCount[26]), 
        .QN(n96) );
  DFFRX1 \inCount_reg[28]  ( .D(N1834), .CK(clk), .RN(n7639), .Q(inCount[28]), 
        .QN(n98) );
  DFFRX1 \inCount_reg[22]  ( .D(N1828), .CK(clk), .RN(n7638), .Q(inCount[22]), 
        .QN(n92) );
  DFFRX1 \inCount_reg[24]  ( .D(N1830), .CK(clk), .RN(n7638), .Q(inCount[24]), 
        .QN(n94) );
  DFFRX1 \inCount_reg[20]  ( .D(N1826), .CK(clk), .RN(n7638), .Q(inCount[20]), 
        .QN(n90) );
  DFFRX1 \inCount_reg[29]  ( .D(N1835), .CK(clk), .RN(n7639), .Q(inCount[29]), 
        .QN(n99) );
  DFFRX1 \inCount_reg[31]  ( .D(N1837), .CK(clk), .RN(n7639), .Q(inCount[31]), 
        .QN(n101) );
  DFFRX1 \inCount_reg[30]  ( .D(N1836), .CK(clk), .RN(n7639), .Q(inCount[30]), 
        .QN(n100) );
  DFFRX1 \inCount_reg[25]  ( .D(N1831), .CK(clk), .RN(n7638), .Q(inCount[25]), 
        .QN(n95) );
  DFFRX1 \inCount_reg[27]  ( .D(N1833), .CK(clk), .RN(n7638), .Q(inCount[27]), 
        .QN(n97) );
  DFFRX1 \inCount_reg[19]  ( .D(N1825), .CK(clk), .RN(n7638), .Q(inCount[19]), 
        .QN(n89) );
  DFFRX1 \inCount_reg[23]  ( .D(N1829), .CK(clk), .RN(n7638), .Q(inCount[23]), 
        .QN(n93) );
  DFFRX1 \outCount_reg[16]  ( .D(outCount_next[16]), .CK(clk), .RN(n7646), .Q(
        outCount[16]) );
  DFFRX1 \outCount_reg[23]  ( .D(outCount_next[23]), .CK(clk), .RN(n7646), .Q(
        outCount[23]) );
  DFFRX1 \outCount_reg[17]  ( .D(outCount_next[17]), .CK(clk), .RN(n7646), .Q(
        outCount[17]) );
  DFFRX1 \outCount_reg[24]  ( .D(outCount_next[24]), .CK(clk), .RN(n7646), .Q(
        outCount[24]) );
  DFFRX1 \outCount_reg[18]  ( .D(outCount_next[18]), .CK(clk), .RN(n7646), .Q(
        outCount[18]) );
  DFFRX1 \outCount_reg[25]  ( .D(outCount_next[25]), .CK(clk), .RN(n7647), .Q(
        outCount[25]) );
  DFFRX1 \outCount_reg[19]  ( .D(outCount_next[19]), .CK(clk), .RN(n7646), .Q(
        outCount[19]) );
  DFFRX1 \outCount_reg[26]  ( .D(outCount_next[26]), .CK(clk), .RN(n7647), .Q(
        outCount[26]) );
  DFFRX1 \outCount_reg[30]  ( .D(outCount_next[30]), .CK(clk), .RN(n7647), .Q(
        outCount[30]) );
  DFFRX1 \outCount_reg[14]  ( .D(outCount_next[14]), .CK(clk), .RN(n7646), .Q(
        outCount[14]) );
  DFFRX1 \outCount_reg[21]  ( .D(outCount_next[21]), .CK(clk), .RN(n7646), .Q(
        outCount[21]) );
  DFFRX1 \outCount_reg[28]  ( .D(outCount_next[28]), .CK(clk), .RN(n7647), .Q(
        outCount[28]) );
  DFFRX1 \outCount_reg[20]  ( .D(outCount_next[20]), .CK(clk), .RN(n7646), .Q(
        outCount[20]) );
  DFFRX1 \outCount_reg[27]  ( .D(outCount_next[27]), .CK(clk), .RN(n7647), .Q(
        outCount[27]) );
  DFFRX1 \outCount_reg[15]  ( .D(outCount_next[15]), .CK(clk), .RN(n7646), .Q(
        outCount[15]) );
  DFFRX1 \outCount_reg[22]  ( .D(outCount_next[22]), .CK(clk), .RN(n7646), .Q(
        outCount[22]) );
  DFFRX1 \outCount_reg[29]  ( .D(outCount_next[29]), .CK(clk), .RN(n7647), .Q(
        outCount[29]) );
  DFFRX1 \state_reg[1]  ( .D(state_next[1]), .CK(clk), .RN(n7639), .Q(state[1]), .QN(n6620) );
  DFFRX1 \state_reg[0]  ( .D(state_next[0]), .CK(clk), .RN(n7639), .Q(state[0]), .QN(n6624) );
  DFFRX1 \xCount_reg[27]  ( .D(xCount_next[27]), .CK(clk), .RN(n7641), .Q(
        xCount[27]), .QN(n130) );
  DFFRX1 \xCount_reg[28]  ( .D(xCount_next[28]), .CK(clk), .RN(n7641), .Q(
        xCount[28]), .QN(n131) );
  DFFRX1 \xCount_reg[22]  ( .D(xCount_next[22]), .CK(clk), .RN(n7641), .Q(
        xCount[22]), .QN(n125) );
  DFFRX1 \xCount_reg[29]  ( .D(xCount_next[29]), .CK(clk), .RN(n7642), .Q(
        xCount[29]), .QN(n132) );
  DFFRX1 \xCount_reg[23]  ( .D(xCount_next[23]), .CK(clk), .RN(n7641), .Q(
        xCount[23]), .QN(n126) );
  DFFRX1 \xCount_reg[30]  ( .D(xCount_next[30]), .CK(clk), .RN(n7642), .Q(
        xCount[30]), .QN(n133) );
  DFFRX1 \iCount_reg[31]  ( .D(n5707), .CK(clk), .RN(n7636), .Q(iCount[31]), 
        .QN(n4902) );
  DFFRX1 \inCount_reg[7]  ( .D(N1813), .CK(clk), .RN(n7637), .Q(inCount[7]), 
        .QN(n77) );
  DFFRX1 \inCount_reg[8]  ( .D(N1814), .CK(clk), .RN(n7637), .Q(inCount[8]), 
        .QN(n78) );
  DFFRX1 \inCount_reg[9]  ( .D(N1815), .CK(clk), .RN(n7637), .Q(inCount[9]), 
        .QN(n79) );
  DFFRX1 \inCount_reg[10]  ( .D(N1816), .CK(clk), .RN(n7637), .Q(inCount[10]), 
        .QN(n80) );
  DFFRX1 \inCount_reg[11]  ( .D(N1817), .CK(clk), .RN(n7637), .Q(inCount[11]), 
        .QN(n81) );
  DFFRX1 \inCount_reg[12]  ( .D(N1818), .CK(clk), .RN(n7637), .Q(inCount[12]), 
        .QN(n82) );
  DFFRX1 \iCount_reg[11]  ( .D(n5727), .CK(clk), .RN(n7634), .Q(iCount[11]), 
        .QN(n4922) );
  DFFRX1 \iCount_reg[14]  ( .D(n5724), .CK(clk), .RN(n7635), .Q(iCount[14]), 
        .QN(n4919) );
  DFFRX1 \iCount_reg[21]  ( .D(n5717), .CK(clk), .RN(n7635), .Q(iCount[21]), 
        .QN(n4912) );
  DFFRX1 \iCount_reg[24]  ( .D(n5714), .CK(clk), .RN(n7636), .Q(iCount[24]), 
        .QN(n4909) );
  DFFRX1 \iCount_reg[27]  ( .D(n5711), .CK(clk), .RN(n7636), .Q(iCount[27]), 
        .QN(n4906) );
  DFFRX1 \outCount_reg[10]  ( .D(outCount_next[10]), .CK(clk), .RN(n7645), .Q(
        outCount[10]) );
  DFFRX1 \iCount_reg[12]  ( .D(n5726), .CK(clk), .RN(n7635), .Q(iCount[12]), 
        .QN(n4921) );
  DFFRX1 \iCount_reg[15]  ( .D(n5723), .CK(clk), .RN(n7635), .Q(iCount[15]), 
        .QN(n4918) );
  DFFRX1 \iCount_reg[22]  ( .D(n5716), .CK(clk), .RN(n7635), .Q(iCount[22]), 
        .QN(n4911) );
  DFFRX1 \iCount_reg[25]  ( .D(n5713), .CK(clk), .RN(n7636), .Q(iCount[25]), 
        .QN(n4908) );
  DFFRX1 \iCount_reg[28]  ( .D(n5710), .CK(clk), .RN(n7636), .Q(iCount[28]), 
        .QN(n4905) );
  DFFRX1 \outCount_reg[11]  ( .D(outCount_next[11]), .CK(clk), .RN(n7645), .Q(
        outCount[11]) );
  DFFRX1 \iCount_reg[13]  ( .D(n5725), .CK(clk), .RN(n7635), .Q(iCount[13]), 
        .QN(n4920) );
  DFFRX1 \iCount_reg[16]  ( .D(n5722), .CK(clk), .RN(n7635), .Q(iCount[16]), 
        .QN(n4917) );
  DFFRX1 \iCount_reg[23]  ( .D(n5715), .CK(clk), .RN(n7635), .Q(iCount[23]), 
        .QN(n4910) );
  DFFRX1 \iCount_reg[26]  ( .D(n5712), .CK(clk), .RN(n7636), .Q(iCount[26]), 
        .QN(n4907) );
  DFFRX1 \iCount_reg[29]  ( .D(n5709), .CK(clk), .RN(n7636), .Q(iCount[29]), 
        .QN(n4904) );
  DFFRX1 \iCount_reg[10]  ( .D(n5728), .CK(clk), .RN(n7634), .Q(iCount[10]), 
        .QN(n4923) );
  DFFRX1 \outCount_reg[12]  ( .D(outCount_next[12]), .CK(clk), .RN(n7645), .Q(
        outCount[12]) );
  DFFRX1 \iCount_reg[17]  ( .D(n5721), .CK(clk), .RN(n7635), .Q(iCount[17]), 
        .QN(n4916) );
  DFFRX1 \iCount_reg[30]  ( .D(n5708), .CK(clk), .RN(n7636), .Q(iCount[30]), 
        .QN(n4903) );
  DFFRX1 \xCount_reg[21]  ( .D(xCount_next[21]), .CK(clk), .RN(n7641), .Q(
        xCount[21]), .QN(n124) );
  DFFRX1 \outCount_reg[8]  ( .D(outCount_next[8]), .CK(clk), .RN(n7645), .Q(
        outCount[8]) );
  DFFRX1 \iCount_reg[8]  ( .D(n5730), .CK(clk), .RN(n7634), .Q(iCount[8]), 
        .QN(n4925) );
  DFFRX1 \iCount_reg[19]  ( .D(n5719), .CK(clk), .RN(n7635), .Q(iCount[19]), 
        .QN(n4914) );
  DFFRX1 \outCount_reg[7]  ( .D(outCount_next[7]), .CK(clk), .RN(n7645), .Q(
        outCount[7]) );
  DFFRX1 \outCount_reg[13]  ( .D(outCount_next[13]), .CK(clk), .RN(n7646), .Q(
        outCount[13]) );
  DFFRX1 \iCount_reg[18]  ( .D(n5720), .CK(clk), .RN(n7635), .Q(iCount[18]), 
        .QN(n4915) );
  DFFRX1 \outCount_reg[9]  ( .D(outCount_next[9]), .CK(clk), .RN(n7645), .Q(
        outCount[9]) );
  DFFRX1 \iCount_reg[9]  ( .D(n5729), .CK(clk), .RN(n7634), .Q(iCount[9]), 
        .QN(n4924) );
  DFFRX1 \iCount_reg[20]  ( .D(n5718), .CK(clk), .RN(n7635), .Q(iCount[20]), 
        .QN(n4913) );
  DFFRX1 doIter_reg ( .D(N1805), .CK(clk), .RN(n7639), .QN(n102) );
  DFFRX1 \xCount_reg[31]  ( .D(xCount_next[31]), .CK(clk), .RN(n7642), .Q(
        xCount[31]) );
  DFFRX1 \xCount_reg[24]  ( .D(xCount_next[24]), .CK(clk), .RN(n7641), .Q(
        xCount[24]) );
  DFFRX1 \inCount_reg[4]  ( .D(N1810), .CK(clk), .RN(n7636), .Q(inCount[4]), 
        .QN(n73) );
  DFFRX1 \inCount_reg[5]  ( .D(N1811), .CK(clk), .RN(n7637), .Q(inCount[5]), 
        .QN(n75) );
  DFFRX1 \inCount_reg[6]  ( .D(N1812), .CK(clk), .RN(n7637), .Q(inCount[6]), 
        .QN(n76) );
  DFFRX1 \iCount_reg[1]  ( .D(n5737), .CK(clk), .RN(n7634), .Q(iCount[1]), 
        .QN(n4932) );
  DFFRX1 \iCount_reg[2]  ( .D(n5736), .CK(clk), .RN(n7634), .Q(iCount[2]), 
        .QN(n4931) );
  DFFRX1 \iCount_reg[3]  ( .D(n5735), .CK(clk), .RN(n7634), .Q(iCount[3]), 
        .QN(n4930) );
  DFFRX1 \iCount_reg[0]  ( .D(n5738), .CK(clk), .RN(n7634), .Q(iCount[0]), 
        .QN(n4933) );
  DFFRX1 \iCount_reg[5]  ( .D(n5733), .CK(clk), .RN(n7634), .Q(iCount[5]), 
        .QN(n4928) );
  DFFRX1 \iCount_reg[4]  ( .D(n5734), .CK(clk), .RN(n7634), .Q(iCount[4]), 
        .QN(n4929) );
  DFFRX1 \outCount_reg[2]  ( .D(outCount_next[2]), .CK(clk), .RN(n7645), .Q(
        outCount[2]) );
  DFFRX1 \outCount_reg[3]  ( .D(outCount_next[3]), .CK(clk), .RN(n7645), .Q(
        outCount[3]) );
  DFFRX1 \outCount_reg[1]  ( .D(n8406), .CK(clk), .RN(n7645), .Q(outCount[1])
         );
  DFFRX1 \xCount_reg[16]  ( .D(xCount_next[16]), .CK(clk), .RN(n7640), .Q(
        xCount[16]), .QN(n119) );
  DFFRX1 \iCount_reg[6]  ( .D(n5732), .CK(clk), .RN(n7634), .Q(iCount[6]), 
        .QN(n4927) );
  DFFRX1 \outCount_reg[6]  ( .D(outCount_next[6]), .CK(clk), .RN(n7645), .Q(
        outCount[6]) );
  DFFRX1 \iCount_reg[7]  ( .D(n5731), .CK(clk), .RN(n7634), .Q(iCount[7]), 
        .QN(n4926) );
  DFFRX1 \outCount_reg[4]  ( .D(outCount_next[4]), .CK(clk), .RN(n7645), .Q(
        outCount[4]) );
  DFFRX1 \xCount_reg[20]  ( .D(xCount_next[20]), .CK(clk), .RN(n7641), .Q(
        xCount[20]), .QN(n123) );
  DFFRX1 \xCount_reg[15]  ( .D(xCount_next[15]), .CK(clk), .RN(n7640), .Q(
        xCount[15]), .QN(n118) );
  DFFRX1 \outCount_reg[5]  ( .D(outCount_next[5]), .CK(clk), .RN(n7645), .Q(
        outCount[5]) );
  DFFRX1 \outCount_reg[0]  ( .D(outCount_next[0]), .CK(clk), .RN(n7644), .Q(
        outCount[0]) );
  DFFRX1 \xCount_reg[17]  ( .D(xCount_next[17]), .CK(clk), .RN(n7641), .Q(
        xCount[17]) );
  DFFRX1 \xCount_reg[19]  ( .D(xCount_next[19]), .CK(clk), .RN(n7641), .Q(
        xCount[19]) );
  DFFRX1 \xCount_reg[26]  ( .D(xCount_next[26]), .CK(clk), .RN(n7641), .Q(
        xCount[26]) );
  DFFRX1 \xCount_reg[18]  ( .D(xCount_next[18]), .CK(clk), .RN(n7641), .Q(
        xCount[18]) );
  DFFRX1 \xCount_reg[25]  ( .D(xCount_next[25]), .CK(clk), .RN(n7641), .Q(
        xCount[25]) );
  DFFRX1 \xCount_reg[8]  ( .D(xCount_next[8]), .CK(clk), .RN(n7640), .Q(
        xCount[8]), .QN(n111) );
  DFFRX1 \xCount_reg[14]  ( .D(xCount_next[14]), .CK(clk), .RN(n7640), .Q(
        xCount[14]), .QN(n117) );
  DFFRX1 \xCount_reg[13]  ( .D(xCount_next[13]), .CK(clk), .RN(n7640), .Q(
        xCount[13]), .QN(n116) );
  DFFRX1 \xCount_reg[9]  ( .D(xCount_next[9]), .CK(clk), .RN(n7640), .Q(
        xCount[9]), .QN(n112) );
  DFFRX1 \xCount_reg[10]  ( .D(xCount_next[10]), .CK(clk), .RN(n7640), .Q(
        xCount[10]) );
  DFFRX1 \xCount_reg[12]  ( .D(xCount_next[12]), .CK(clk), .RN(n7640), .Q(
        xCount[12]) );
  DFFRX1 \xCount_reg[11]  ( .D(xCount_next[11]), .CK(clk), .RN(n7640), .Q(
        xCount[11]) );
  DFFRX1 \xCount_reg[6]  ( .D(xCount_next[6]), .CK(clk), .RN(n7640), .Q(
        xCount[6]), .QN(n109) );
  DFFRX1 \xCount_reg[7]  ( .D(xCount_next[7]), .CK(clk), .RN(n7640), .Q(
        xCount[7]), .QN(n110) );
  DFFRX1 \xCount_reg[5]  ( .D(xCount_next[5]), .CK(clk), .RN(n7640), .Q(
        xCount[5]) );
  DFFRX1 \xCount_reg[4]  ( .D(xCount_next[4]), .CK(clk), .RN(n7639), .Q(
        xCount[4]) );
  DFFQX1 \xArray_reg[1][63]  ( .D(N28768), .CK(clk), .Q(\xArray[1][63] ) );
  DFFQX1 \xArray_reg[13][63]  ( .D(N28000), .CK(clk), .Q(\xArray[13][63] ) );
  DFFQX1 \xArray_reg[9][63]  ( .D(N28256), .CK(clk), .Q(\xArray[9][63] ) );
  DFFQX1 \xArray_reg[8][63]  ( .D(N28320), .CK(clk), .Q(\xArray[8][63] ) );
  DFFRX1 \bArray_reg[1][63]  ( .D(n6458), .CK(clk), .RN(n7574), .Q(
        \bArray[1][63] ), .QN(n5653) );
  DFFRX1 \bArray_reg[1][62]  ( .D(n6457), .CK(clk), .RN(n7574), .Q(
        \bArray[1][62] ), .QN(n5652) );
  DFFRX1 \bArray_reg[1][61]  ( .D(n6456), .CK(clk), .RN(n7574), .Q(
        \bArray[1][61] ), .QN(n5651) );
  DFFRX1 \bArray_reg[1][60]  ( .D(n6455), .CK(clk), .RN(n7574), .Q(
        \bArray[1][60] ), .QN(n5650) );
  DFFRX1 \bArray_reg[5][63]  ( .D(n6266), .CK(clk), .RN(n7590), .Q(
        \bArray[5][63] ), .QN(n5461) );
  DFFRX1 \bArray_reg[5][62]  ( .D(n6265), .CK(clk), .RN(n7590), .Q(
        \bArray[5][62] ), .QN(n5460) );
  DFFRX1 \bArray_reg[5][61]  ( .D(n6264), .CK(clk), .RN(n7590), .Q(
        \bArray[5][61] ), .QN(n5459) );
  DFFRX1 \bArray_reg[5][60]  ( .D(n6263), .CK(clk), .RN(n7590), .Q(
        \bArray[5][60] ), .QN(n5458) );
  DFFRX1 \bArray_reg[9][63]  ( .D(n6074), .CK(clk), .RN(n7606), .Q(
        \bArray[9][63] ), .QN(n5269) );
  DFFRX1 \bArray_reg[9][62]  ( .D(n6073), .CK(clk), .RN(n7606), .Q(
        \bArray[9][62] ), .QN(n5268) );
  DFFRX1 \bArray_reg[9][61]  ( .D(n6072), .CK(clk), .RN(n7606), .Q(
        \bArray[9][61] ), .QN(n5267) );
  DFFRX1 \bArray_reg[9][60]  ( .D(n6071), .CK(clk), .RN(n7606), .Q(
        \bArray[9][60] ), .QN(n5266) );
  DFFRX1 \bArray_reg[13][63]  ( .D(n5882), .CK(clk), .RN(n7622), .Q(
        \bArray[13][63] ), .QN(n5077) );
  DFFRX1 \bArray_reg[13][62]  ( .D(n5881), .CK(clk), .RN(n7622), .Q(
        \bArray[13][62] ), .QN(n5076) );
  DFFRX1 \bArray_reg[13][61]  ( .D(n5880), .CK(clk), .RN(n7622), .Q(
        \bArray[13][61] ), .QN(n5075) );
  DFFRX1 \bArray_reg[13][60]  ( .D(n5879), .CK(clk), .RN(n7622), .Q(
        \bArray[13][60] ), .QN(n5074) );
  DFFRX1 \bArray_reg[3][63]  ( .D(n6362), .CK(clk), .RN(n7582), .Q(
        \bArray[3][63] ), .QN(n5557) );
  DFFRX1 \bArray_reg[3][62]  ( .D(n6361), .CK(clk), .RN(n7582), .Q(
        \bArray[3][62] ), .QN(n5556) );
  DFFRX1 \bArray_reg[3][61]  ( .D(n6360), .CK(clk), .RN(n7582), .Q(
        \bArray[3][61] ), .QN(n5555) );
  DFFRX1 \bArray_reg[3][60]  ( .D(n6359), .CK(clk), .RN(n7582), .Q(
        \bArray[3][60] ), .QN(n5554) );
  DFFRX1 \bArray_reg[7][63]  ( .D(n6170), .CK(clk), .RN(n7598), .Q(
        \bArray[7][63] ), .QN(n5365) );
  DFFRX1 \bArray_reg[7][62]  ( .D(n6169), .CK(clk), .RN(n7598), .Q(
        \bArray[7][62] ), .QN(n5364) );
  DFFRX1 \bArray_reg[7][61]  ( .D(n6168), .CK(clk), .RN(n7598), .Q(
        \bArray[7][61] ), .QN(n5363) );
  DFFRX1 \bArray_reg[7][60]  ( .D(n6167), .CK(clk), .RN(n7598), .Q(
        \bArray[7][60] ), .QN(n5362) );
  DFFRX1 \bArray_reg[11][63]  ( .D(n5978), .CK(clk), .RN(n7614), .Q(
        \bArray[11][63] ), .QN(n5173) );
  DFFRX1 \bArray_reg[11][62]  ( .D(n5977), .CK(clk), .RN(n7614), .Q(
        \bArray[11][62] ), .QN(n5172) );
  DFFRX1 \bArray_reg[11][61]  ( .D(n5976), .CK(clk), .RN(n7614), .Q(
        \bArray[11][61] ), .QN(n5171) );
  DFFRX1 \bArray_reg[11][60]  ( .D(n5975), .CK(clk), .RN(n7614), .Q(
        \bArray[11][60] ), .QN(n5170) );
  DFFRX1 \bArray_reg[15][63]  ( .D(n5786), .CK(clk), .RN(n7630), .Q(
        \bArray[15][63] ), .QN(n4981) );
  DFFRX1 \bArray_reg[15][62]  ( .D(n5785), .CK(clk), .RN(n7630), .Q(
        \bArray[15][62] ), .QN(n4980) );
  DFFRX1 \bArray_reg[15][61]  ( .D(n5784), .CK(clk), .RN(n7630), .Q(
        \bArray[15][61] ), .QN(n4979) );
  DFFRX1 \bArray_reg[15][60]  ( .D(n5783), .CK(clk), .RN(n7630), .Q(
        \bArray[15][60] ), .QN(n4978) );
  DFFRX1 \bArray_reg[0][63]  ( .D(n6506), .CK(clk), .RN(n7570), .Q(
        \bArray[0][63] ), .QN(n5704) );
  DFFRX1 \bArray_reg[0][62]  ( .D(n6505), .CK(clk), .RN(n7570), .Q(
        \bArray[0][62] ), .QN(n5700) );
  DFFRX1 \bArray_reg[0][61]  ( .D(n6504), .CK(clk), .RN(n7570), .Q(
        \bArray[0][61] ), .QN(n5699) );
  DFFRX1 \bArray_reg[0][60]  ( .D(n6503), .CK(clk), .RN(n7570), .Q(
        \bArray[0][60] ), .QN(n5698) );
  DFFRX1 \bArray_reg[4][63]  ( .D(n6314), .CK(clk), .RN(n7586), .Q(
        \bArray[4][63] ), .QN(n5509) );
  DFFRX1 \bArray_reg[4][62]  ( .D(n6313), .CK(clk), .RN(n7586), .Q(
        \bArray[4][62] ), .QN(n5508) );
  DFFRX1 \bArray_reg[4][61]  ( .D(n6312), .CK(clk), .RN(n7586), .Q(
        \bArray[4][61] ), .QN(n5507) );
  DFFRX1 \bArray_reg[4][60]  ( .D(n6311), .CK(clk), .RN(n7586), .Q(
        \bArray[4][60] ), .QN(n5506) );
  DFFRX1 \bArray_reg[8][63]  ( .D(n6122), .CK(clk), .RN(n7602), .Q(
        \bArray[8][63] ), .QN(n5317) );
  DFFRX1 \bArray_reg[8][62]  ( .D(n6121), .CK(clk), .RN(n7602), .Q(
        \bArray[8][62] ), .QN(n5316) );
  DFFRX1 \bArray_reg[8][61]  ( .D(n6120), .CK(clk), .RN(n7602), .Q(
        \bArray[8][61] ), .QN(n5315) );
  DFFRX1 \bArray_reg[8][60]  ( .D(n6119), .CK(clk), .RN(n7602), .Q(
        \bArray[8][60] ), .QN(n5314) );
  DFFRX1 \bArray_reg[12][63]  ( .D(n5930), .CK(clk), .RN(n7618), .Q(
        \bArray[12][63] ), .QN(n5125) );
  DFFRX1 \bArray_reg[12][62]  ( .D(n5929), .CK(clk), .RN(n7618), .Q(
        \bArray[12][62] ), .QN(n5124) );
  DFFRX1 \bArray_reg[12][61]  ( .D(n5928), .CK(clk), .RN(n7618), .Q(
        \bArray[12][61] ), .QN(n5123) );
  DFFRX1 \bArray_reg[12][60]  ( .D(n5927), .CK(clk), .RN(n7618), .Q(
        \bArray[12][60] ), .QN(n5122) );
  DFFRX1 \bArray_reg[2][63]  ( .D(n6410), .CK(clk), .RN(n7578), .Q(
        \bArray[2][63] ), .QN(n5605) );
  DFFRX1 \bArray_reg[2][62]  ( .D(n6409), .CK(clk), .RN(n7578), .Q(
        \bArray[2][62] ), .QN(n5604) );
  DFFRX1 \bArray_reg[2][61]  ( .D(n6408), .CK(clk), .RN(n7578), .Q(
        \bArray[2][61] ), .QN(n5603) );
  DFFRX1 \bArray_reg[2][60]  ( .D(n6407), .CK(clk), .RN(n7578), .Q(
        \bArray[2][60] ), .QN(n5602) );
  DFFRX1 \bArray_reg[6][63]  ( .D(n6218), .CK(clk), .RN(n7594), .Q(
        \bArray[6][63] ), .QN(n5413) );
  DFFRX1 \bArray_reg[6][62]  ( .D(n6217), .CK(clk), .RN(n7594), .Q(
        \bArray[6][62] ), .QN(n5412) );
  DFFRX1 \bArray_reg[6][61]  ( .D(n6216), .CK(clk), .RN(n7594), .Q(
        \bArray[6][61] ), .QN(n5411) );
  DFFRX1 \bArray_reg[10][63]  ( .D(n6026), .CK(clk), .RN(n7610), .Q(
        \bArray[10][63] ), .QN(n5221) );
  DFFRX1 \bArray_reg[10][62]  ( .D(n6025), .CK(clk), .RN(n7610), .Q(
        \bArray[10][62] ), .QN(n5220) );
  DFFRX1 \bArray_reg[10][61]  ( .D(n6024), .CK(clk), .RN(n7610), .Q(
        \bArray[10][61] ), .QN(n5219) );
  DFFRX1 \bArray_reg[10][60]  ( .D(n6023), .CK(clk), .RN(n7610), .Q(
        \bArray[10][60] ), .QN(n5218) );
  DFFRX1 \bArray_reg[14][63]  ( .D(n5834), .CK(clk), .RN(n7626), .Q(
        \bArray[14][63] ), .QN(n5029) );
  DFFRX1 \bArray_reg[14][62]  ( .D(n5833), .CK(clk), .RN(n7626), .Q(
        \bArray[14][62] ), .QN(n5028) );
  DFFRX1 \bArray_reg[14][61]  ( .D(n5832), .CK(clk), .RN(n7626), .Q(
        \bArray[14][61] ), .QN(n5027) );
  DFFRX1 \bArray_reg[14][60]  ( .D(n5831), .CK(clk), .RN(n7626), .Q(
        \bArray[14][60] ), .QN(n5026) );
  DFFRX1 \bArray_reg[6][60]  ( .D(n6215), .CK(clk), .RN(n7594), .Q(
        \bArray[6][60] ), .QN(n5410) );
  DFFQX1 \xArray_reg[1][62]  ( .D(N28767), .CK(clk), .Q(\xArray[1][62] ) );
  DFFQX1 \xArray_reg[13][62]  ( .D(N27999), .CK(clk), .Q(\xArray[13][62] ) );
  DFFQX1 \xArray_reg[9][62]  ( .D(N28255), .CK(clk), .Q(\xArray[9][62] ) );
  DFFQX1 \xArray_reg[8][62]  ( .D(N28319), .CK(clk), .Q(\xArray[8][62] ) );
  DFFRX1 \bArray_reg[1][59]  ( .D(n6454), .CK(clk), .RN(n7574), .Q(
        \bArray[1][59] ), .QN(n5649) );
  DFFRX1 \bArray_reg[1][58]  ( .D(n6453), .CK(clk), .RN(n7574), .Q(
        \bArray[1][58] ), .QN(n5648) );
  DFFRX1 \bArray_reg[1][57]  ( .D(n6452), .CK(clk), .RN(n7574), .Q(
        \bArray[1][57] ), .QN(n5647) );
  DFFRX1 \bArray_reg[1][56]  ( .D(n6451), .CK(clk), .RN(n7574), .Q(
        \bArray[1][56] ), .QN(n5646) );
  DFFRX1 \bArray_reg[5][59]  ( .D(n6262), .CK(clk), .RN(n7590), .Q(
        \bArray[5][59] ), .QN(n5457) );
  DFFRX1 \bArray_reg[5][58]  ( .D(n6261), .CK(clk), .RN(n7590), .Q(
        \bArray[5][58] ), .QN(n5456) );
  DFFRX1 \bArray_reg[5][57]  ( .D(n6260), .CK(clk), .RN(n7590), .Q(
        \bArray[5][57] ), .QN(n5455) );
  DFFRX1 \bArray_reg[5][56]  ( .D(n6259), .CK(clk), .RN(n7590), .Q(
        \bArray[5][56] ), .QN(n5454) );
  DFFRX1 \bArray_reg[9][59]  ( .D(n6070), .CK(clk), .RN(n7606), .Q(
        \bArray[9][59] ), .QN(n5265) );
  DFFRX1 \bArray_reg[9][58]  ( .D(n6069), .CK(clk), .RN(n7606), .Q(
        \bArray[9][58] ), .QN(n5264) );
  DFFRX1 \bArray_reg[9][57]  ( .D(n6068), .CK(clk), .RN(n7606), .Q(
        \bArray[9][57] ), .QN(n5263) );
  DFFRX1 \bArray_reg[9][56]  ( .D(n6067), .CK(clk), .RN(n7606), .Q(
        \bArray[9][56] ), .QN(n5262) );
  DFFRX1 \bArray_reg[13][59]  ( .D(n5878), .CK(clk), .RN(n7622), .Q(
        \bArray[13][59] ), .QN(n5073) );
  DFFRX1 \bArray_reg[13][58]  ( .D(n5877), .CK(clk), .RN(n7622), .Q(
        \bArray[13][58] ), .QN(n5072) );
  DFFRX1 \bArray_reg[13][57]  ( .D(n5876), .CK(clk), .RN(n7622), .Q(
        \bArray[13][57] ), .QN(n5071) );
  DFFRX1 \bArray_reg[13][56]  ( .D(n5875), .CK(clk), .RN(n7622), .Q(
        \bArray[13][56] ), .QN(n5070) );
  DFFRX1 \bArray_reg[3][59]  ( .D(n6358), .CK(clk), .RN(n7582), .Q(
        \bArray[3][59] ), .QN(n5553) );
  DFFRX1 \bArray_reg[3][58]  ( .D(n6357), .CK(clk), .RN(n7582), .Q(
        \bArray[3][58] ), .QN(n5552) );
  DFFRX1 \bArray_reg[3][57]  ( .D(n6356), .CK(clk), .RN(n7582), .Q(
        \bArray[3][57] ), .QN(n5551) );
  DFFRX1 \bArray_reg[3][56]  ( .D(n6355), .CK(clk), .RN(n7582), .Q(
        \bArray[3][56] ), .QN(n5550) );
  DFFRX1 \bArray_reg[7][59]  ( .D(n6166), .CK(clk), .RN(n7598), .Q(
        \bArray[7][59] ), .QN(n5361) );
  DFFRX1 \bArray_reg[7][58]  ( .D(n6165), .CK(clk), .RN(n7598), .Q(
        \bArray[7][58] ), .QN(n5360) );
  DFFRX1 \bArray_reg[7][57]  ( .D(n6164), .CK(clk), .RN(n7598), .Q(
        \bArray[7][57] ), .QN(n5359) );
  DFFRX1 \bArray_reg[7][56]  ( .D(n6163), .CK(clk), .RN(n7598), .Q(
        \bArray[7][56] ), .QN(n5358) );
  DFFRX1 \bArray_reg[11][59]  ( .D(n5974), .CK(clk), .RN(n7614), .Q(
        \bArray[11][59] ), .QN(n5169) );
  DFFRX1 \bArray_reg[11][58]  ( .D(n5973), .CK(clk), .RN(n7614), .Q(
        \bArray[11][58] ), .QN(n5168) );
  DFFRX1 \bArray_reg[11][57]  ( .D(n5972), .CK(clk), .RN(n7614), .Q(
        \bArray[11][57] ), .QN(n5167) );
  DFFRX1 \bArray_reg[11][56]  ( .D(n5971), .CK(clk), .RN(n7614), .Q(
        \bArray[11][56] ), .QN(n5166) );
  DFFRX1 \bArray_reg[15][59]  ( .D(n5782), .CK(clk), .RN(n7630), .Q(
        \bArray[15][59] ), .QN(n4977) );
  DFFRX1 \bArray_reg[15][58]  ( .D(n5781), .CK(clk), .RN(n7630), .Q(
        \bArray[15][58] ), .QN(n4976) );
  DFFRX1 \bArray_reg[15][57]  ( .D(n5780), .CK(clk), .RN(n7630), .Q(
        \bArray[15][57] ), .QN(n4975) );
  DFFRX1 \bArray_reg[15][56]  ( .D(n5779), .CK(clk), .RN(n7630), .Q(
        \bArray[15][56] ), .QN(n4974) );
  DFFRX1 \bArray_reg[0][59]  ( .D(n6502), .CK(clk), .RN(n7570), .Q(
        \bArray[0][59] ), .QN(n5697) );
  DFFRX1 \bArray_reg[0][58]  ( .D(n6501), .CK(clk), .RN(n7570), .Q(
        \bArray[0][58] ), .QN(n5696) );
  DFFRX1 \bArray_reg[0][57]  ( .D(n6500), .CK(clk), .RN(n7570), .Q(
        \bArray[0][57] ), .QN(n5695) );
  DFFRX1 \bArray_reg[0][56]  ( .D(n6499), .CK(clk), .RN(n7570), .Q(
        \bArray[0][56] ), .QN(n5694) );
  DFFRX1 \bArray_reg[4][59]  ( .D(n6310), .CK(clk), .RN(n7586), .Q(
        \bArray[4][59] ), .QN(n5505) );
  DFFRX1 \bArray_reg[4][58]  ( .D(n6309), .CK(clk), .RN(n7586), .Q(
        \bArray[4][58] ), .QN(n5504) );
  DFFRX1 \bArray_reg[4][57]  ( .D(n6308), .CK(clk), .RN(n7586), .Q(
        \bArray[4][57] ), .QN(n5503) );
  DFFRX1 \bArray_reg[4][56]  ( .D(n6307), .CK(clk), .RN(n7586), .Q(
        \bArray[4][56] ), .QN(n5502) );
  DFFRX1 \bArray_reg[8][59]  ( .D(n6118), .CK(clk), .RN(n7602), .Q(
        \bArray[8][59] ), .QN(n5313) );
  DFFRX1 \bArray_reg[8][58]  ( .D(n6117), .CK(clk), .RN(n7602), .Q(
        \bArray[8][58] ), .QN(n5312) );
  DFFRX1 \bArray_reg[8][57]  ( .D(n6116), .CK(clk), .RN(n7602), .Q(
        \bArray[8][57] ), .QN(n5311) );
  DFFRX1 \bArray_reg[8][56]  ( .D(n6115), .CK(clk), .RN(n7602), .Q(
        \bArray[8][56] ), .QN(n5310) );
  DFFRX1 \bArray_reg[12][59]  ( .D(n5926), .CK(clk), .RN(n7618), .Q(
        \bArray[12][59] ), .QN(n5121) );
  DFFRX1 \bArray_reg[12][58]  ( .D(n5925), .CK(clk), .RN(n7618), .Q(
        \bArray[12][58] ), .QN(n5120) );
  DFFRX1 \bArray_reg[12][57]  ( .D(n5924), .CK(clk), .RN(n7618), .Q(
        \bArray[12][57] ), .QN(n5119) );
  DFFRX1 \bArray_reg[12][56]  ( .D(n5923), .CK(clk), .RN(n7618), .Q(
        \bArray[12][56] ), .QN(n5118) );
  DFFRX1 \bArray_reg[2][59]  ( .D(n6406), .CK(clk), .RN(n7578), .Q(
        \bArray[2][59] ), .QN(n5601) );
  DFFRX1 \bArray_reg[2][58]  ( .D(n6405), .CK(clk), .RN(n7578), .Q(
        \bArray[2][58] ), .QN(n5600) );
  DFFRX1 \bArray_reg[2][57]  ( .D(n6404), .CK(clk), .RN(n7578), .Q(
        \bArray[2][57] ), .QN(n5599) );
  DFFRX1 \bArray_reg[2][56]  ( .D(n6403), .CK(clk), .RN(n7578), .Q(
        \bArray[2][56] ), .QN(n5598) );
  DFFRX1 \bArray_reg[6][59]  ( .D(n6214), .CK(clk), .RN(n7594), .Q(
        \bArray[6][59] ), .QN(n5409) );
  DFFRX1 \bArray_reg[6][58]  ( .D(n6213), .CK(clk), .RN(n7594), .Q(
        \bArray[6][58] ), .QN(n5408) );
  DFFRX1 \bArray_reg[6][57]  ( .D(n6212), .CK(clk), .RN(n7594), .Q(
        \bArray[6][57] ), .QN(n5407) );
  DFFRX1 \bArray_reg[6][56]  ( .D(n6211), .CK(clk), .RN(n7594), .Q(
        \bArray[6][56] ), .QN(n5406) );
  DFFRX1 \bArray_reg[10][59]  ( .D(n6022), .CK(clk), .RN(n7610), .Q(
        \bArray[10][59] ), .QN(n5217) );
  DFFRX1 \bArray_reg[10][58]  ( .D(n6021), .CK(clk), .RN(n7610), .Q(
        \bArray[10][58] ), .QN(n5216) );
  DFFRX1 \bArray_reg[10][57]  ( .D(n6020), .CK(clk), .RN(n7610), .Q(
        \bArray[10][57] ), .QN(n5215) );
  DFFRX1 \bArray_reg[10][56]  ( .D(n6019), .CK(clk), .RN(n7610), .Q(
        \bArray[10][56] ), .QN(n5214) );
  DFFRX1 \bArray_reg[14][59]  ( .D(n5830), .CK(clk), .RN(n7626), .Q(
        \bArray[14][59] ), .QN(n5025) );
  DFFRX1 \bArray_reg[14][58]  ( .D(n5829), .CK(clk), .RN(n7626), .Q(
        \bArray[14][58] ), .QN(n5024) );
  DFFRX1 \bArray_reg[14][57]  ( .D(n5828), .CK(clk), .RN(n7626), .Q(
        \bArray[14][57] ), .QN(n5023) );
  DFFRX1 \bArray_reg[14][56]  ( .D(n5827), .CK(clk), .RN(n7626), .Q(
        \bArray[14][56] ), .QN(n5022) );
  DFFQX1 \xArray_reg[1][61]  ( .D(N28766), .CK(clk), .Q(\xArray[1][61] ) );
  DFFQX1 \xArray_reg[13][61]  ( .D(N27998), .CK(clk), .Q(\xArray[13][61] ) );
  DFFQX1 \xArray_reg[9][61]  ( .D(N28254), .CK(clk), .Q(\xArray[9][61] ) );
  DFFQX1 \xArray_reg[8][61]  ( .D(N28318), .CK(clk), .Q(\xArray[8][61] ) );
  DFFQX1 \xArray_reg[9][60]  ( .D(N28253), .CK(clk), .Q(\xArray[9][60] ) );
  DFFQX1 \xArray_reg[8][60]  ( .D(N28317), .CK(clk), .Q(\xArray[8][60] ) );
  DFFRX1 \bArray_reg[1][55]  ( .D(n6450), .CK(clk), .RN(n7574), .Q(
        \bArray[1][55] ), .QN(n5645) );
  DFFRX1 \bArray_reg[1][54]  ( .D(n6449), .CK(clk), .RN(n7574), .Q(
        \bArray[1][54] ), .QN(n5644) );
  DFFRX1 \bArray_reg[1][53]  ( .D(n6448), .CK(clk), .RN(n7574), .Q(
        \bArray[1][53] ), .QN(n5643) );
  DFFRX1 \bArray_reg[1][52]  ( .D(n6447), .CK(clk), .RN(n7574), .Q(
        \bArray[1][52] ), .QN(n5642) );
  DFFRX1 \bArray_reg[5][55]  ( .D(n6258), .CK(clk), .RN(n7590), .Q(
        \bArray[5][55] ), .QN(n5453) );
  DFFRX1 \bArray_reg[5][54]  ( .D(n6257), .CK(clk), .RN(n7590), .Q(
        \bArray[5][54] ), .QN(n5452) );
  DFFRX1 \bArray_reg[5][53]  ( .D(n6256), .CK(clk), .RN(n7590), .Q(
        \bArray[5][53] ), .QN(n5451) );
  DFFRX1 \bArray_reg[5][52]  ( .D(n6255), .CK(clk), .RN(n7590), .Q(
        \bArray[5][52] ), .QN(n5450) );
  DFFRX1 \bArray_reg[9][55]  ( .D(n6066), .CK(clk), .RN(n7606), .Q(
        \bArray[9][55] ), .QN(n5261) );
  DFFRX1 \bArray_reg[9][54]  ( .D(n6065), .CK(clk), .RN(n7606), .Q(
        \bArray[9][54] ), .QN(n5260) );
  DFFRX1 \bArray_reg[9][53]  ( .D(n6064), .CK(clk), .RN(n7606), .Q(
        \bArray[9][53] ), .QN(n5259) );
  DFFRX1 \bArray_reg[9][52]  ( .D(n6063), .CK(clk), .RN(n7606), .Q(
        \bArray[9][52] ), .QN(n5258) );
  DFFRX1 \bArray_reg[13][55]  ( .D(n5874), .CK(clk), .RN(n7622), .Q(
        \bArray[13][55] ), .QN(n5069) );
  DFFRX1 \bArray_reg[13][54]  ( .D(n5873), .CK(clk), .RN(n7622), .Q(
        \bArray[13][54] ), .QN(n5068) );
  DFFRX1 \bArray_reg[13][53]  ( .D(n5872), .CK(clk), .RN(n7622), .Q(
        \bArray[13][53] ), .QN(n5067) );
  DFFRX1 \bArray_reg[13][52]  ( .D(n5871), .CK(clk), .RN(n7622), .Q(
        \bArray[13][52] ), .QN(n5066) );
  DFFRX1 \bArray_reg[3][55]  ( .D(n6354), .CK(clk), .RN(n7582), .Q(
        \bArray[3][55] ), .QN(n5549) );
  DFFRX1 \bArray_reg[3][54]  ( .D(n6353), .CK(clk), .RN(n7582), .Q(
        \bArray[3][54] ), .QN(n5548) );
  DFFRX1 \bArray_reg[3][53]  ( .D(n6352), .CK(clk), .RN(n7582), .Q(
        \bArray[3][53] ), .QN(n5547) );
  DFFRX1 \bArray_reg[3][52]  ( .D(n6351), .CK(clk), .RN(n7582), .Q(
        \bArray[3][52] ), .QN(n5546) );
  DFFRX1 \bArray_reg[7][55]  ( .D(n6162), .CK(clk), .RN(n7598), .Q(
        \bArray[7][55] ), .QN(n5357) );
  DFFRX1 \bArray_reg[7][54]  ( .D(n6161), .CK(clk), .RN(n7598), .Q(
        \bArray[7][54] ), .QN(n5356) );
  DFFRX1 \bArray_reg[7][53]  ( .D(n6160), .CK(clk), .RN(n7598), .Q(
        \bArray[7][53] ), .QN(n5355) );
  DFFRX1 \bArray_reg[7][52]  ( .D(n6159), .CK(clk), .RN(n7598), .Q(
        \bArray[7][52] ), .QN(n5354) );
  DFFRX1 \bArray_reg[11][55]  ( .D(n5970), .CK(clk), .RN(n7614), .Q(
        \bArray[11][55] ), .QN(n5165) );
  DFFRX1 \bArray_reg[11][54]  ( .D(n5969), .CK(clk), .RN(n7614), .Q(
        \bArray[11][54] ), .QN(n5164) );
  DFFRX1 \bArray_reg[11][53]  ( .D(n5968), .CK(clk), .RN(n7614), .Q(
        \bArray[11][53] ), .QN(n5163) );
  DFFRX1 \bArray_reg[11][52]  ( .D(n5967), .CK(clk), .RN(n7614), .Q(
        \bArray[11][52] ), .QN(n5162) );
  DFFRX1 \bArray_reg[15][55]  ( .D(n5778), .CK(clk), .RN(n7630), .Q(
        \bArray[15][55] ), .QN(n4973) );
  DFFRX1 \bArray_reg[15][54]  ( .D(n5777), .CK(clk), .RN(n7630), .Q(
        \bArray[15][54] ), .QN(n4972) );
  DFFRX1 \bArray_reg[15][53]  ( .D(n5776), .CK(clk), .RN(n7630), .Q(
        \bArray[15][53] ), .QN(n4971) );
  DFFRX1 \bArray_reg[15][52]  ( .D(n5775), .CK(clk), .RN(n7630), .Q(
        \bArray[15][52] ), .QN(n4970) );
  DFFRX1 \bArray_reg[0][55]  ( .D(n6498), .CK(clk), .RN(n7570), .Q(
        \bArray[0][55] ), .QN(n5693) );
  DFFRX1 \bArray_reg[0][54]  ( .D(n6497), .CK(clk), .RN(n7570), .Q(
        \bArray[0][54] ), .QN(n5692) );
  DFFRX1 \bArray_reg[0][53]  ( .D(n6496), .CK(clk), .RN(n7570), .Q(
        \bArray[0][53] ), .QN(n5691) );
  DFFRX1 \bArray_reg[0][52]  ( .D(n6495), .CK(clk), .RN(n7570), .Q(
        \bArray[0][52] ), .QN(n5690) );
  DFFRX1 \bArray_reg[4][55]  ( .D(n6306), .CK(clk), .RN(n7586), .Q(
        \bArray[4][55] ), .QN(n5501) );
  DFFRX1 \bArray_reg[4][54]  ( .D(n6305), .CK(clk), .RN(n7586), .Q(
        \bArray[4][54] ), .QN(n5500) );
  DFFRX1 \bArray_reg[4][53]  ( .D(n6304), .CK(clk), .RN(n7586), .Q(
        \bArray[4][53] ), .QN(n5499) );
  DFFRX1 \bArray_reg[4][52]  ( .D(n6303), .CK(clk), .RN(n7586), .Q(
        \bArray[4][52] ), .QN(n5498) );
  DFFRX1 \bArray_reg[8][55]  ( .D(n6114), .CK(clk), .RN(n7602), .Q(
        \bArray[8][55] ), .QN(n5309) );
  DFFRX1 \bArray_reg[8][54]  ( .D(n6113), .CK(clk), .RN(n7602), .Q(
        \bArray[8][54] ), .QN(n5308) );
  DFFRX1 \bArray_reg[8][53]  ( .D(n6112), .CK(clk), .RN(n7602), .Q(
        \bArray[8][53] ), .QN(n5307) );
  DFFRX1 \bArray_reg[8][52]  ( .D(n6111), .CK(clk), .RN(n7602), .Q(
        \bArray[8][52] ), .QN(n5306) );
  DFFRX1 \bArray_reg[12][55]  ( .D(n5922), .CK(clk), .RN(n7618), .Q(
        \bArray[12][55] ), .QN(n5117) );
  DFFRX1 \bArray_reg[12][54]  ( .D(n5921), .CK(clk), .RN(n7618), .Q(
        \bArray[12][54] ), .QN(n5116) );
  DFFRX1 \bArray_reg[12][53]  ( .D(n5920), .CK(clk), .RN(n7618), .Q(
        \bArray[12][53] ), .QN(n5115) );
  DFFRX1 \bArray_reg[12][52]  ( .D(n5919), .CK(clk), .RN(n7618), .Q(
        \bArray[12][52] ), .QN(n5114) );
  DFFRX1 \bArray_reg[2][55]  ( .D(n6402), .CK(clk), .RN(n7578), .Q(
        \bArray[2][55] ), .QN(n5597) );
  DFFRX1 \bArray_reg[2][54]  ( .D(n6401), .CK(clk), .RN(n7578), .Q(
        \bArray[2][54] ), .QN(n5596) );
  DFFRX1 \bArray_reg[2][53]  ( .D(n6400), .CK(clk), .RN(n7578), .Q(
        \bArray[2][53] ), .QN(n5595) );
  DFFRX1 \bArray_reg[2][52]  ( .D(n6399), .CK(clk), .RN(n7578), .Q(
        \bArray[2][52] ), .QN(n5594) );
  DFFRX1 \bArray_reg[6][55]  ( .D(n6210), .CK(clk), .RN(n7594), .Q(
        \bArray[6][55] ), .QN(n5405) );
  DFFRX1 \bArray_reg[6][54]  ( .D(n6209), .CK(clk), .RN(n7594), .Q(
        \bArray[6][54] ), .QN(n5404) );
  DFFRX1 \bArray_reg[6][53]  ( .D(n6208), .CK(clk), .RN(n7594), .Q(
        \bArray[6][53] ), .QN(n5403) );
  DFFRX1 \bArray_reg[6][52]  ( .D(n6207), .CK(clk), .RN(n7594), .Q(
        \bArray[6][52] ), .QN(n5402) );
  DFFRX1 \bArray_reg[10][55]  ( .D(n6018), .CK(clk), .RN(n7610), .Q(
        \bArray[10][55] ), .QN(n5213) );
  DFFRX1 \bArray_reg[10][54]  ( .D(n6017), .CK(clk), .RN(n7610), .Q(
        \bArray[10][54] ), .QN(n5212) );
  DFFRX1 \bArray_reg[10][53]  ( .D(n6016), .CK(clk), .RN(n7610), .Q(
        \bArray[10][53] ), .QN(n5211) );
  DFFRX1 \bArray_reg[10][52]  ( .D(n6015), .CK(clk), .RN(n7610), .Q(
        \bArray[10][52] ), .QN(n5210) );
  DFFRX1 \bArray_reg[14][55]  ( .D(n5826), .CK(clk), .RN(n7626), .Q(
        \bArray[14][55] ), .QN(n5021) );
  DFFRX1 \bArray_reg[14][54]  ( .D(n5825), .CK(clk), .RN(n7626), .Q(
        \bArray[14][54] ), .QN(n5020) );
  DFFRX1 \bArray_reg[14][53]  ( .D(n5824), .CK(clk), .RN(n7626), .Q(
        \bArray[14][53] ), .QN(n5019) );
  DFFRX1 \bArray_reg[14][52]  ( .D(n5823), .CK(clk), .RN(n7626), .Q(
        \bArray[14][52] ), .QN(n5018) );
  DFFQX1 \xArray_reg[1][60]  ( .D(N28765), .CK(clk), .Q(\xArray[1][60] ) );
  DFFQX1 \xArray_reg[1][59]  ( .D(N28764), .CK(clk), .Q(\xArray[1][59] ) );
  DFFQX1 \xArray_reg[13][60]  ( .D(N27997), .CK(clk), .Q(\xArray[13][60] ) );
  DFFQX1 \xArray_reg[13][59]  ( .D(N27996), .CK(clk), .Q(\xArray[13][59] ) );
  DFFQX1 \xArray_reg[9][59]  ( .D(N28252), .CK(clk), .Q(\xArray[9][59] ) );
  DFFQX1 \xArray_reg[9][58]  ( .D(N28251), .CK(clk), .Q(\xArray[9][58] ) );
  DFFQX1 \xArray_reg[8][59]  ( .D(N28316), .CK(clk), .Q(\xArray[8][59] ) );
  DFFQX1 \xArray_reg[8][58]  ( .D(N28315), .CK(clk), .Q(\xArray[8][58] ) );
  DFFQX1 \xArray_reg[1][58]  ( .D(N28763), .CK(clk), .Q(\xArray[1][58] ) );
  DFFQX1 \xArray_reg[1][57]  ( .D(N28762), .CK(clk), .Q(\xArray[1][57] ) );
  DFFQX1 \xArray_reg[13][58]  ( .D(N27995), .CK(clk), .Q(\xArray[13][58] ) );
  DFFQX1 \xArray_reg[13][57]  ( .D(N27994), .CK(clk), .Q(\xArray[13][57] ) );
  DFFQX1 \xArray_reg[9][57]  ( .D(N28250), .CK(clk), .Q(\xArray[9][57] ) );
  DFFQX1 \xArray_reg[9][56]  ( .D(N28249), .CK(clk), .Q(\xArray[9][56] ) );
  DFFQX1 \xArray_reg[8][57]  ( .D(N28314), .CK(clk), .Q(\xArray[8][57] ) );
  DFFQX1 \xArray_reg[8][56]  ( .D(N28313), .CK(clk), .Q(\xArray[8][56] ) );
  DFFRX1 \bArray_reg[1][51]  ( .D(n6446), .CK(clk), .RN(n7575), .Q(
        \bArray[1][51] ), .QN(n5641) );
  DFFRX1 \bArray_reg[1][50]  ( .D(n6445), .CK(clk), .RN(n7575), .Q(
        \bArray[1][50] ), .QN(n5640) );
  DFFRX1 \bArray_reg[1][49]  ( .D(n6444), .CK(clk), .RN(n7575), .Q(
        \bArray[1][49] ), .QN(n5639) );
  DFFRX1 \bArray_reg[1][48]  ( .D(n6443), .CK(clk), .RN(n7575), .Q(
        \bArray[1][48] ), .QN(n5638) );
  DFFRX1 \bArray_reg[5][51]  ( .D(n6254), .CK(clk), .RN(n7591), .Q(
        \bArray[5][51] ), .QN(n5449) );
  DFFRX1 \bArray_reg[5][50]  ( .D(n6253), .CK(clk), .RN(n7591), .Q(
        \bArray[5][50] ), .QN(n5448) );
  DFFRX1 \bArray_reg[5][49]  ( .D(n6252), .CK(clk), .RN(n7591), .Q(
        \bArray[5][49] ), .QN(n5447) );
  DFFRX1 \bArray_reg[5][48]  ( .D(n6251), .CK(clk), .RN(n7591), .Q(
        \bArray[5][48] ), .QN(n5446) );
  DFFRX1 \bArray_reg[9][51]  ( .D(n6062), .CK(clk), .RN(n7607), .Q(
        \bArray[9][51] ), .QN(n5257) );
  DFFRX1 \bArray_reg[9][50]  ( .D(n6061), .CK(clk), .RN(n7607), .Q(
        \bArray[9][50] ), .QN(n5256) );
  DFFRX1 \bArray_reg[9][49]  ( .D(n6060), .CK(clk), .RN(n7607), .Q(
        \bArray[9][49] ), .QN(n5255) );
  DFFRX1 \bArray_reg[9][48]  ( .D(n6059), .CK(clk), .RN(n7607), .Q(
        \bArray[9][48] ), .QN(n5254) );
  DFFRX1 \bArray_reg[13][51]  ( .D(n5870), .CK(clk), .RN(n7623), .Q(
        \bArray[13][51] ), .QN(n5065) );
  DFFRX1 \bArray_reg[13][50]  ( .D(n5869), .CK(clk), .RN(n7623), .Q(
        \bArray[13][50] ), .QN(n5064) );
  DFFRX1 \bArray_reg[13][49]  ( .D(n5868), .CK(clk), .RN(n7623), .Q(
        \bArray[13][49] ), .QN(n5063) );
  DFFRX1 \bArray_reg[13][48]  ( .D(n5867), .CK(clk), .RN(n7623), .Q(
        \bArray[13][48] ), .QN(n5062) );
  DFFRX1 \bArray_reg[3][51]  ( .D(n6350), .CK(clk), .RN(n7583), .Q(
        \bArray[3][51] ), .QN(n5545) );
  DFFRX1 \bArray_reg[3][50]  ( .D(n6349), .CK(clk), .RN(n7583), .Q(
        \bArray[3][50] ), .QN(n5544) );
  DFFRX1 \bArray_reg[3][49]  ( .D(n6348), .CK(clk), .RN(n7583), .Q(
        \bArray[3][49] ), .QN(n5543) );
  DFFRX1 \bArray_reg[3][48]  ( .D(n6347), .CK(clk), .RN(n7583), .Q(
        \bArray[3][48] ), .QN(n5542) );
  DFFRX1 \bArray_reg[7][51]  ( .D(n6158), .CK(clk), .RN(n7599), .Q(
        \bArray[7][51] ), .QN(n5353) );
  DFFRX1 \bArray_reg[7][50]  ( .D(n6157), .CK(clk), .RN(n7599), .Q(
        \bArray[7][50] ), .QN(n5352) );
  DFFRX1 \bArray_reg[7][49]  ( .D(n6156), .CK(clk), .RN(n7599), .Q(
        \bArray[7][49] ), .QN(n5351) );
  DFFRX1 \bArray_reg[7][48]  ( .D(n6155), .CK(clk), .RN(n7599), .Q(
        \bArray[7][48] ), .QN(n5350) );
  DFFRX1 \bArray_reg[11][51]  ( .D(n5966), .CK(clk), .RN(n7615), .Q(
        \bArray[11][51] ), .QN(n5161) );
  DFFRX1 \bArray_reg[11][50]  ( .D(n5965), .CK(clk), .RN(n7615), .Q(
        \bArray[11][50] ), .QN(n5160) );
  DFFRX1 \bArray_reg[11][49]  ( .D(n5964), .CK(clk), .RN(n7615), .Q(
        \bArray[11][49] ), .QN(n5159) );
  DFFRX1 \bArray_reg[11][48]  ( .D(n5963), .CK(clk), .RN(n7615), .Q(
        \bArray[11][48] ), .QN(n5158) );
  DFFRX1 \bArray_reg[15][51]  ( .D(n5774), .CK(clk), .RN(n7631), .Q(
        \bArray[15][51] ), .QN(n4969) );
  DFFRX1 \bArray_reg[15][50]  ( .D(n5773), .CK(clk), .RN(n7631), .Q(
        \bArray[15][50] ), .QN(n4968) );
  DFFRX1 \bArray_reg[15][49]  ( .D(n5772), .CK(clk), .RN(n7631), .Q(
        \bArray[15][49] ), .QN(n4967) );
  DFFRX1 \bArray_reg[15][48]  ( .D(n5771), .CK(clk), .RN(n7631), .Q(
        \bArray[15][48] ), .QN(n4966) );
  DFFRX1 \bArray_reg[0][51]  ( .D(n6494), .CK(clk), .RN(n7571), .Q(
        \bArray[0][51] ), .QN(n5689) );
  DFFRX1 \bArray_reg[0][50]  ( .D(n6493), .CK(clk), .RN(n7571), .Q(
        \bArray[0][50] ), .QN(n5688) );
  DFFRX1 \bArray_reg[0][49]  ( .D(n6492), .CK(clk), .RN(n7571), .Q(
        \bArray[0][49] ), .QN(n5687) );
  DFFRX1 \bArray_reg[0][48]  ( .D(n6491), .CK(clk), .RN(n7571), .Q(
        \bArray[0][48] ), .QN(n5686) );
  DFFRX1 \bArray_reg[4][51]  ( .D(n6302), .CK(clk), .RN(n7587), .Q(
        \bArray[4][51] ), .QN(n5497) );
  DFFRX1 \bArray_reg[4][50]  ( .D(n6301), .CK(clk), .RN(n7587), .Q(
        \bArray[4][50] ), .QN(n5496) );
  DFFRX1 \bArray_reg[4][49]  ( .D(n6300), .CK(clk), .RN(n7587), .Q(
        \bArray[4][49] ), .QN(n5495) );
  DFFRX1 \bArray_reg[4][48]  ( .D(n6299), .CK(clk), .RN(n7587), .Q(
        \bArray[4][48] ), .QN(n5494) );
  DFFRX1 \bArray_reg[8][51]  ( .D(n6110), .CK(clk), .RN(n7603), .Q(
        \bArray[8][51] ), .QN(n5305) );
  DFFRX1 \bArray_reg[8][50]  ( .D(n6109), .CK(clk), .RN(n7603), .Q(
        \bArray[8][50] ), .QN(n5304) );
  DFFRX1 \bArray_reg[8][49]  ( .D(n6108), .CK(clk), .RN(n7603), .Q(
        \bArray[8][49] ), .QN(n5303) );
  DFFRX1 \bArray_reg[8][48]  ( .D(n6107), .CK(clk), .RN(n7603), .Q(
        \bArray[8][48] ), .QN(n5302) );
  DFFRX1 \bArray_reg[12][51]  ( .D(n5918), .CK(clk), .RN(n7619), .Q(
        \bArray[12][51] ), .QN(n5113) );
  DFFRX1 \bArray_reg[12][50]  ( .D(n5917), .CK(clk), .RN(n7619), .Q(
        \bArray[12][50] ), .QN(n5112) );
  DFFRX1 \bArray_reg[12][49]  ( .D(n5916), .CK(clk), .RN(n7619), .Q(
        \bArray[12][49] ), .QN(n5111) );
  DFFRX1 \bArray_reg[12][48]  ( .D(n5915), .CK(clk), .RN(n7619), .Q(
        \bArray[12][48] ), .QN(n5110) );
  DFFRX1 \bArray_reg[2][51]  ( .D(n6398), .CK(clk), .RN(n7579), .Q(
        \bArray[2][51] ), .QN(n5593) );
  DFFRX1 \bArray_reg[2][50]  ( .D(n6397), .CK(clk), .RN(n7579), .Q(
        \bArray[2][50] ), .QN(n5592) );
  DFFRX1 \bArray_reg[2][49]  ( .D(n6396), .CK(clk), .RN(n7579), .Q(
        \bArray[2][49] ), .QN(n5591) );
  DFFRX1 \bArray_reg[2][48]  ( .D(n6395), .CK(clk), .RN(n7579), .Q(
        \bArray[2][48] ), .QN(n5590) );
  DFFRX1 \bArray_reg[6][51]  ( .D(n6206), .CK(clk), .RN(n7595), .Q(
        \bArray[6][51] ), .QN(n5401) );
  DFFRX1 \bArray_reg[6][50]  ( .D(n6205), .CK(clk), .RN(n7595), .Q(
        \bArray[6][50] ), .QN(n5400) );
  DFFRX1 \bArray_reg[6][49]  ( .D(n6204), .CK(clk), .RN(n7595), .Q(
        \bArray[6][49] ), .QN(n5399) );
  DFFRX1 \bArray_reg[6][48]  ( .D(n6203), .CK(clk), .RN(n7595), .Q(
        \bArray[6][48] ), .QN(n5398) );
  DFFRX1 \bArray_reg[10][51]  ( .D(n6014), .CK(clk), .RN(n7611), .Q(
        \bArray[10][51] ), .QN(n5209) );
  DFFRX1 \bArray_reg[10][50]  ( .D(n6013), .CK(clk), .RN(n7611), .Q(
        \bArray[10][50] ), .QN(n5208) );
  DFFRX1 \bArray_reg[10][49]  ( .D(n6012), .CK(clk), .RN(n7611), .Q(
        \bArray[10][49] ), .QN(n5207) );
  DFFRX1 \bArray_reg[10][48]  ( .D(n6011), .CK(clk), .RN(n7611), .Q(
        \bArray[10][48] ), .QN(n5206) );
  DFFRX1 \bArray_reg[14][51]  ( .D(n5822), .CK(clk), .RN(n7627), .Q(
        \bArray[14][51] ), .QN(n5017) );
  DFFRX1 \bArray_reg[14][50]  ( .D(n5821), .CK(clk), .RN(n7627), .Q(
        \bArray[14][50] ), .QN(n5016) );
  DFFRX1 \bArray_reg[14][49]  ( .D(n5820), .CK(clk), .RN(n7627), .Q(
        \bArray[14][49] ), .QN(n5015) );
  DFFRX1 \bArray_reg[14][48]  ( .D(n5819), .CK(clk), .RN(n7627), .Q(
        \bArray[14][48] ), .QN(n5014) );
  DFFQX1 \xArray_reg[1][56]  ( .D(N28761), .CK(clk), .Q(\xArray[1][56] ) );
  DFFQX1 \xArray_reg[1][55]  ( .D(N28760), .CK(clk), .Q(\xArray[1][55] ) );
  DFFQX1 \xArray_reg[1][54]  ( .D(N28759), .CK(clk), .Q(\xArray[1][54] ) );
  DFFQX1 \xArray_reg[13][56]  ( .D(N27993), .CK(clk), .Q(\xArray[13][56] ) );
  DFFQX1 \xArray_reg[13][55]  ( .D(N27992), .CK(clk), .Q(\xArray[13][55] ) );
  DFFQX1 \xArray_reg[13][54]  ( .D(N27991), .CK(clk), .Q(\xArray[13][54] ) );
  DFFQX1 \xArray_reg[9][55]  ( .D(N28248), .CK(clk), .Q(\xArray[9][55] ) );
  DFFQX1 \xArray_reg[9][54]  ( .D(N28247), .CK(clk), .Q(\xArray[9][54] ) );
  DFFQX1 \xArray_reg[9][53]  ( .D(N28246), .CK(clk), .Q(\xArray[9][53] ) );
  DFFQX1 \xArray_reg[8][55]  ( .D(N28312), .CK(clk), .Q(\xArray[8][55] ) );
  DFFQX1 \xArray_reg[8][54]  ( .D(N28311), .CK(clk), .Q(\xArray[8][54] ) );
  DFFQX1 \xArray_reg[8][53]  ( .D(N28310), .CK(clk), .Q(\xArray[8][53] ) );
  DFFQX1 \xArray_reg[1][53]  ( .D(N28758), .CK(clk), .Q(\xArray[1][53] ) );
  DFFQX1 \xArray_reg[1][52]  ( .D(N28757), .CK(clk), .Q(\xArray[1][52] ) );
  DFFQX1 \xArray_reg[13][53]  ( .D(N27990), .CK(clk), .Q(\xArray[13][53] ) );
  DFFQX1 \xArray_reg[13][52]  ( .D(N27989), .CK(clk), .Q(\xArray[13][52] ) );
  DFFQX1 \xArray_reg[9][52]  ( .D(N28245), .CK(clk), .Q(\xArray[9][52] ) );
  DFFQX1 \xArray_reg[8][52]  ( .D(N28309), .CK(clk), .Q(\xArray[8][52] ) );
  DFFRX1 \bArray_reg[1][47]  ( .D(n6442), .CK(clk), .RN(n7575), .Q(
        \bArray[1][47] ), .QN(n5637) );
  DFFRX1 \bArray_reg[1][46]  ( .D(n6441), .CK(clk), .RN(n7575), .Q(
        \bArray[1][46] ), .QN(n5636) );
  DFFRX1 \bArray_reg[1][45]  ( .D(n6440), .CK(clk), .RN(n7575), .Q(
        \bArray[1][45] ), .QN(n5635) );
  DFFRX1 \bArray_reg[1][44]  ( .D(n6439), .CK(clk), .RN(n7575), .Q(
        \bArray[1][44] ), .QN(n5634) );
  DFFRX1 \bArray_reg[5][47]  ( .D(n6250), .CK(clk), .RN(n7591), .Q(
        \bArray[5][47] ), .QN(n5445) );
  DFFRX1 \bArray_reg[5][46]  ( .D(n6249), .CK(clk), .RN(n7591), .Q(
        \bArray[5][46] ), .QN(n5444) );
  DFFRX1 \bArray_reg[5][45]  ( .D(n6248), .CK(clk), .RN(n7591), .Q(
        \bArray[5][45] ), .QN(n5443) );
  DFFRX1 \bArray_reg[5][44]  ( .D(n6247), .CK(clk), .RN(n7591), .Q(
        \bArray[5][44] ), .QN(n5442) );
  DFFRX1 \bArray_reg[9][47]  ( .D(n6058), .CK(clk), .RN(n7607), .Q(
        \bArray[9][47] ), .QN(n5253) );
  DFFRX1 \bArray_reg[9][46]  ( .D(n6057), .CK(clk), .RN(n7607), .Q(
        \bArray[9][46] ), .QN(n5252) );
  DFFRX1 \bArray_reg[9][45]  ( .D(n6056), .CK(clk), .RN(n7607), .Q(
        \bArray[9][45] ), .QN(n5251) );
  DFFRX1 \bArray_reg[9][44]  ( .D(n6055), .CK(clk), .RN(n7607), .Q(
        \bArray[9][44] ), .QN(n5250) );
  DFFRX1 \bArray_reg[13][47]  ( .D(n5866), .CK(clk), .RN(n7623), .Q(
        \bArray[13][47] ), .QN(n5061) );
  DFFRX1 \bArray_reg[13][46]  ( .D(n5865), .CK(clk), .RN(n7623), .Q(
        \bArray[13][46] ), .QN(n5060) );
  DFFRX1 \bArray_reg[13][45]  ( .D(n5864), .CK(clk), .RN(n7623), .Q(
        \bArray[13][45] ), .QN(n5059) );
  DFFRX1 \bArray_reg[13][44]  ( .D(n5863), .CK(clk), .RN(n7623), .Q(
        \bArray[13][44] ), .QN(n5058) );
  DFFRX1 \bArray_reg[3][47]  ( .D(n6346), .CK(clk), .RN(n7583), .Q(
        \bArray[3][47] ), .QN(n5541) );
  DFFRX1 \bArray_reg[3][46]  ( .D(n6345), .CK(clk), .RN(n7583), .Q(
        \bArray[3][46] ), .QN(n5540) );
  DFFRX1 \bArray_reg[3][45]  ( .D(n6344), .CK(clk), .RN(n7583), .Q(
        \bArray[3][45] ), .QN(n5539) );
  DFFRX1 \bArray_reg[3][44]  ( .D(n6343), .CK(clk), .RN(n7583), .Q(
        \bArray[3][44] ), .QN(n5538) );
  DFFRX1 \bArray_reg[7][47]  ( .D(n6154), .CK(clk), .RN(n7599), .Q(
        \bArray[7][47] ), .QN(n5349) );
  DFFRX1 \bArray_reg[7][46]  ( .D(n6153), .CK(clk), .RN(n7599), .Q(
        \bArray[7][46] ), .QN(n5348) );
  DFFRX1 \bArray_reg[7][45]  ( .D(n6152), .CK(clk), .RN(n7599), .Q(
        \bArray[7][45] ), .QN(n5347) );
  DFFRX1 \bArray_reg[7][44]  ( .D(n6151), .CK(clk), .RN(n7599), .Q(
        \bArray[7][44] ), .QN(n5346) );
  DFFRX1 \bArray_reg[11][47]  ( .D(n5962), .CK(clk), .RN(n7615), .Q(
        \bArray[11][47] ), .QN(n5157) );
  DFFRX1 \bArray_reg[11][46]  ( .D(n5961), .CK(clk), .RN(n7615), .Q(
        \bArray[11][46] ), .QN(n5156) );
  DFFRX1 \bArray_reg[11][45]  ( .D(n5960), .CK(clk), .RN(n7615), .Q(
        \bArray[11][45] ), .QN(n5155) );
  DFFRX1 \bArray_reg[11][44]  ( .D(n5959), .CK(clk), .RN(n7615), .Q(
        \bArray[11][44] ), .QN(n5154) );
  DFFRX1 \bArray_reg[15][47]  ( .D(n5770), .CK(clk), .RN(n7631), .Q(
        \bArray[15][47] ), .QN(n4965) );
  DFFRX1 \bArray_reg[15][46]  ( .D(n5769), .CK(clk), .RN(n7631), .Q(
        \bArray[15][46] ), .QN(n4964) );
  DFFRX1 \bArray_reg[15][45]  ( .D(n5768), .CK(clk), .RN(n7631), .Q(
        \bArray[15][45] ), .QN(n4963) );
  DFFRX1 \bArray_reg[15][44]  ( .D(n5767), .CK(clk), .RN(n7631), .Q(
        \bArray[15][44] ), .QN(n4962) );
  DFFRX1 \bArray_reg[0][47]  ( .D(n6490), .CK(clk), .RN(n7571), .Q(
        \bArray[0][47] ), .QN(n5685) );
  DFFRX1 \bArray_reg[0][46]  ( .D(n6489), .CK(clk), .RN(n7571), .Q(
        \bArray[0][46] ), .QN(n5684) );
  DFFRX1 \bArray_reg[0][45]  ( .D(n6488), .CK(clk), .RN(n7571), .Q(
        \bArray[0][45] ), .QN(n5683) );
  DFFRX1 \bArray_reg[0][44]  ( .D(n6487), .CK(clk), .RN(n7571), .Q(
        \bArray[0][44] ), .QN(n5682) );
  DFFRX1 \bArray_reg[4][47]  ( .D(n6298), .CK(clk), .RN(n7587), .Q(
        \bArray[4][47] ), .QN(n5493) );
  DFFRX1 \bArray_reg[4][46]  ( .D(n6297), .CK(clk), .RN(n7587), .Q(
        \bArray[4][46] ), .QN(n5492) );
  DFFRX1 \bArray_reg[4][45]  ( .D(n6296), .CK(clk), .RN(n7587), .Q(
        \bArray[4][45] ), .QN(n5491) );
  DFFRX1 \bArray_reg[4][44]  ( .D(n6295), .CK(clk), .RN(n7587), .Q(
        \bArray[4][44] ), .QN(n5490) );
  DFFRX1 \bArray_reg[8][47]  ( .D(n6106), .CK(clk), .RN(n7603), .Q(
        \bArray[8][47] ), .QN(n5301) );
  DFFRX1 \bArray_reg[8][46]  ( .D(n6105), .CK(clk), .RN(n7603), .Q(
        \bArray[8][46] ), .QN(n5300) );
  DFFRX1 \bArray_reg[8][45]  ( .D(n6104), .CK(clk), .RN(n7603), .Q(
        \bArray[8][45] ), .QN(n5299) );
  DFFRX1 \bArray_reg[8][44]  ( .D(n6103), .CK(clk), .RN(n7603), .Q(
        \bArray[8][44] ), .QN(n5298) );
  DFFRX1 \bArray_reg[12][47]  ( .D(n5914), .CK(clk), .RN(n7619), .Q(
        \bArray[12][47] ), .QN(n5109) );
  DFFRX1 \bArray_reg[12][46]  ( .D(n5913), .CK(clk), .RN(n7619), .Q(
        \bArray[12][46] ), .QN(n5108) );
  DFFRX1 \bArray_reg[12][45]  ( .D(n5912), .CK(clk), .RN(n7619), .Q(
        \bArray[12][45] ), .QN(n5107) );
  DFFRX1 \bArray_reg[12][44]  ( .D(n5911), .CK(clk), .RN(n7619), .Q(
        \bArray[12][44] ), .QN(n5106) );
  DFFRX1 \bArray_reg[2][47]  ( .D(n6394), .CK(clk), .RN(n7579), .Q(
        \bArray[2][47] ), .QN(n5589) );
  DFFRX1 \bArray_reg[2][46]  ( .D(n6393), .CK(clk), .RN(n7579), .Q(
        \bArray[2][46] ), .QN(n5588) );
  DFFRX1 \bArray_reg[2][45]  ( .D(n6392), .CK(clk), .RN(n7579), .Q(
        \bArray[2][45] ), .QN(n5587) );
  DFFRX1 \bArray_reg[2][44]  ( .D(n6391), .CK(clk), .RN(n7579), .Q(
        \bArray[2][44] ), .QN(n5586) );
  DFFRX1 \bArray_reg[6][47]  ( .D(n6202), .CK(clk), .RN(n7595), .Q(
        \bArray[6][47] ), .QN(n5397) );
  DFFRX1 \bArray_reg[6][46]  ( .D(n6201), .CK(clk), .RN(n7595), .Q(
        \bArray[6][46] ), .QN(n5396) );
  DFFRX1 \bArray_reg[6][45]  ( .D(n6200), .CK(clk), .RN(n7595), .Q(
        \bArray[6][45] ), .QN(n5395) );
  DFFRX1 \bArray_reg[6][44]  ( .D(n6199), .CK(clk), .RN(n7595), .Q(
        \bArray[6][44] ), .QN(n5394) );
  DFFRX1 \bArray_reg[10][47]  ( .D(n6010), .CK(clk), .RN(n7611), .Q(
        \bArray[10][47] ), .QN(n5205) );
  DFFRX1 \bArray_reg[10][46]  ( .D(n6009), .CK(clk), .RN(n7611), .Q(
        \bArray[10][46] ), .QN(n5204) );
  DFFRX1 \bArray_reg[10][45]  ( .D(n6008), .CK(clk), .RN(n7611), .Q(
        \bArray[10][45] ), .QN(n5203) );
  DFFRX1 \bArray_reg[10][44]  ( .D(n6007), .CK(clk), .RN(n7611), .Q(
        \bArray[10][44] ), .QN(n5202) );
  DFFRX1 \bArray_reg[14][47]  ( .D(n5818), .CK(clk), .RN(n7627), .Q(
        \bArray[14][47] ), .QN(n5013) );
  DFFRX1 \bArray_reg[14][46]  ( .D(n5817), .CK(clk), .RN(n7627), .Q(
        \bArray[14][46] ), .QN(n5012) );
  DFFRX1 \bArray_reg[14][45]  ( .D(n5816), .CK(clk), .RN(n7627), .Q(
        \bArray[14][45] ), .QN(n5011) );
  DFFRX1 \bArray_reg[14][44]  ( .D(n5815), .CK(clk), .RN(n7627), .Q(
        \bArray[14][44] ), .QN(n5010) );
  DFFQX1 \xArray_reg[1][51]  ( .D(N28756), .CK(clk), .Q(\xArray[1][51] ) );
  DFFQX1 \xArray_reg[1][50]  ( .D(N28755), .CK(clk), .Q(\xArray[1][50] ) );
  DFFQX1 \xArray_reg[13][51]  ( .D(N27988), .CK(clk), .Q(\xArray[13][51] ) );
  DFFQX1 \xArray_reg[13][50]  ( .D(N27987), .CK(clk), .Q(\xArray[13][50] ) );
  DFFQX1 \xArray_reg[9][51]  ( .D(N28244), .CK(clk), .Q(\xArray[9][51] ) );
  DFFQX1 \xArray_reg[9][50]  ( .D(N28243), .CK(clk), .Q(\xArray[9][50] ) );
  DFFQX1 \xArray_reg[8][51]  ( .D(N28308), .CK(clk), .Q(\xArray[8][51] ) );
  DFFQX1 \xArray_reg[8][50]  ( .D(N28307), .CK(clk), .Q(\xArray[8][50] ) );
  DFFQX1 \xArray_reg[3][48]  ( .D(N28625), .CK(clk), .Q(\xArray[3][48] ) );
  DFFQX1 \xArray_reg[3][47]  ( .D(N28624), .CK(clk), .Q(\xArray[3][47] ) );
  DFFQX1 \xArray_reg[15][48]  ( .D(N27857), .CK(clk), .Q(\xArray[15][48] ) );
  DFFQX1 \xArray_reg[0][48]  ( .D(N28817), .CK(clk), .Q(\xArray[0][48] ) );
  DFFQX1 \xArray_reg[4][48]  ( .D(N28561), .CK(clk), .Q(\xArray[4][48] ) );
  DFFQX1 \xArray_reg[5][48]  ( .D(N28497), .CK(clk), .Q(\xArray[5][48] ) );
  DFFQX1 \xArray_reg[14][48]  ( .D(N27921), .CK(clk), .Q(\xArray[14][48] ) );
  DFFQX1 \xArray_reg[11][48]  ( .D(N28113), .CK(clk), .Q(\xArray[11][48] ) );
  DFFQX1 \xArray_reg[12][48]  ( .D(N28049), .CK(clk), .Q(\xArray[12][48] ) );
  DFFQX1 \xArray_reg[7][48]  ( .D(N28369), .CK(clk), .Q(\xArray[7][48] ) );
  DFFQX1 \xArray_reg[7][47]  ( .D(N28368), .CK(clk), .Q(\xArray[7][47] ) );
  DFFQX1 \xArray_reg[1][49]  ( .D(N28754), .CK(clk), .Q(\xArray[1][49] ) );
  DFFQX1 \xArray_reg[1][48]  ( .D(N28753), .CK(clk), .Q(\xArray[1][48] ) );
  DFFQX1 \xArray_reg[13][49]  ( .D(N27986), .CK(clk), .Q(\xArray[13][49] ) );
  DFFQX1 \xArray_reg[13][48]  ( .D(N27985), .CK(clk), .Q(\xArray[13][48] ) );
  DFFQX1 \xArray_reg[9][49]  ( .D(N28242), .CK(clk), .Q(\xArray[9][49] ) );
  DFFQX1 \xArray_reg[9][48]  ( .D(N28241), .CK(clk), .Q(\xArray[9][48] ) );
  DFFQX1 \xArray_reg[8][49]  ( .D(N28306), .CK(clk), .Q(\xArray[8][49] ) );
  DFFQX1 \xArray_reg[8][48]  ( .D(N28305), .CK(clk), .Q(\xArray[8][48] ) );
  DFFQX1 \xArray_reg[10][48]  ( .D(N28177), .CK(clk), .Q(\xArray[10][48] ) );
  DFFQX1 \xArray_reg[10][47]  ( .D(N28176), .CK(clk), .Q(\xArray[10][47] ) );
  DFFQX1 \xArray_reg[6][48]  ( .D(N28433), .CK(clk), .Q(\xArray[6][48] ) );
  DFFQX1 \xArray_reg[6][47]  ( .D(N28432), .CK(clk), .Q(\xArray[6][47] ) );
  DFFRX1 \bArray_reg[1][43]  ( .D(n6438), .CK(clk), .RN(n7575), .Q(
        \bArray[1][43] ), .QN(n5633) );
  DFFRX1 \bArray_reg[1][42]  ( .D(n6437), .CK(clk), .RN(n7575), .Q(
        \bArray[1][42] ), .QN(n5632) );
  DFFRX1 \bArray_reg[1][41]  ( .D(n6436), .CK(clk), .RN(n7575), .Q(
        \bArray[1][41] ), .QN(n5631) );
  DFFRX1 \bArray_reg[1][40]  ( .D(n6435), .CK(clk), .RN(n7575), .Q(
        \bArray[1][40] ), .QN(n5630) );
  DFFRX1 \bArray_reg[5][43]  ( .D(n6246), .CK(clk), .RN(n7591), .Q(
        \bArray[5][43] ), .QN(n5441) );
  DFFRX1 \bArray_reg[5][42]  ( .D(n6245), .CK(clk), .RN(n7591), .Q(
        \bArray[5][42] ), .QN(n5440) );
  DFFRX1 \bArray_reg[5][41]  ( .D(n6244), .CK(clk), .RN(n7591), .Q(
        \bArray[5][41] ), .QN(n5439) );
  DFFRX1 \bArray_reg[5][40]  ( .D(n6243), .CK(clk), .RN(n7591), .Q(
        \bArray[5][40] ), .QN(n5438) );
  DFFRX1 \bArray_reg[9][43]  ( .D(n6054), .CK(clk), .RN(n7607), .Q(
        \bArray[9][43] ), .QN(n5249) );
  DFFRX1 \bArray_reg[9][42]  ( .D(n6053), .CK(clk), .RN(n7607), .Q(
        \bArray[9][42] ), .QN(n5248) );
  DFFRX1 \bArray_reg[9][41]  ( .D(n6052), .CK(clk), .RN(n7607), .Q(
        \bArray[9][41] ), .QN(n5247) );
  DFFRX1 \bArray_reg[9][40]  ( .D(n6051), .CK(clk), .RN(n7607), .Q(
        \bArray[9][40] ), .QN(n5246) );
  DFFRX1 \bArray_reg[13][43]  ( .D(n5862), .CK(clk), .RN(n7623), .Q(
        \bArray[13][43] ), .QN(n5057) );
  DFFRX1 \bArray_reg[13][42]  ( .D(n5861), .CK(clk), .RN(n7623), .Q(
        \bArray[13][42] ), .QN(n5056) );
  DFFRX1 \bArray_reg[13][41]  ( .D(n5860), .CK(clk), .RN(n7623), .Q(
        \bArray[13][41] ), .QN(n5055) );
  DFFRX1 \bArray_reg[13][40]  ( .D(n5859), .CK(clk), .RN(n7623), .Q(
        \bArray[13][40] ), .QN(n5054) );
  DFFRX1 \bArray_reg[3][43]  ( .D(n6342), .CK(clk), .RN(n7583), .Q(
        \bArray[3][43] ), .QN(n5537) );
  DFFRX1 \bArray_reg[3][42]  ( .D(n6341), .CK(clk), .RN(n7583), .Q(
        \bArray[3][42] ), .QN(n5536) );
  DFFRX1 \bArray_reg[3][41]  ( .D(n6340), .CK(clk), .RN(n7583), .Q(
        \bArray[3][41] ), .QN(n5535) );
  DFFRX1 \bArray_reg[3][40]  ( .D(n6339), .CK(clk), .RN(n7583), .Q(
        \bArray[3][40] ), .QN(n5534) );
  DFFRX1 \bArray_reg[7][43]  ( .D(n6150), .CK(clk), .RN(n7599), .Q(
        \bArray[7][43] ), .QN(n5345) );
  DFFRX1 \bArray_reg[7][42]  ( .D(n6149), .CK(clk), .RN(n7599), .Q(
        \bArray[7][42] ), .QN(n5344) );
  DFFRX1 \bArray_reg[7][41]  ( .D(n6148), .CK(clk), .RN(n7599), .Q(
        \bArray[7][41] ), .QN(n5343) );
  DFFRX1 \bArray_reg[7][40]  ( .D(n6147), .CK(clk), .RN(n7599), .Q(
        \bArray[7][40] ), .QN(n5342) );
  DFFRX1 \bArray_reg[11][43]  ( .D(n5958), .CK(clk), .RN(n7615), .Q(
        \bArray[11][43] ), .QN(n5153) );
  DFFRX1 \bArray_reg[11][42]  ( .D(n5957), .CK(clk), .RN(n7615), .Q(
        \bArray[11][42] ), .QN(n5152) );
  DFFRX1 \bArray_reg[11][41]  ( .D(n5956), .CK(clk), .RN(n7615), .Q(
        \bArray[11][41] ), .QN(n5151) );
  DFFRX1 \bArray_reg[11][40]  ( .D(n5955), .CK(clk), .RN(n7615), .Q(
        \bArray[11][40] ), .QN(n5150) );
  DFFRX1 \bArray_reg[15][43]  ( .D(n5766), .CK(clk), .RN(n7631), .Q(
        \bArray[15][43] ), .QN(n4961) );
  DFFRX1 \bArray_reg[15][42]  ( .D(n5765), .CK(clk), .RN(n7631), .Q(
        \bArray[15][42] ), .QN(n4960) );
  DFFRX1 \bArray_reg[15][41]  ( .D(n5764), .CK(clk), .RN(n7631), .Q(
        \bArray[15][41] ), .QN(n4959) );
  DFFRX1 \bArray_reg[15][40]  ( .D(n5763), .CK(clk), .RN(n7631), .Q(
        \bArray[15][40] ), .QN(n4958) );
  DFFRX1 \bArray_reg[0][43]  ( .D(n6486), .CK(clk), .RN(n7571), .Q(
        \bArray[0][43] ), .QN(n5681) );
  DFFRX1 \bArray_reg[0][42]  ( .D(n6485), .CK(clk), .RN(n7571), .Q(
        \bArray[0][42] ), .QN(n5680) );
  DFFRX1 \bArray_reg[0][41]  ( .D(n6484), .CK(clk), .RN(n7571), .Q(
        \bArray[0][41] ), .QN(n5679) );
  DFFRX1 \bArray_reg[0][40]  ( .D(n6483), .CK(clk), .RN(n7571), .Q(
        \bArray[0][40] ), .QN(n5678) );
  DFFRX1 \bArray_reg[4][43]  ( .D(n6294), .CK(clk), .RN(n7587), .Q(
        \bArray[4][43] ), .QN(n5489) );
  DFFRX1 \bArray_reg[4][42]  ( .D(n6293), .CK(clk), .RN(n7587), .Q(
        \bArray[4][42] ), .QN(n5488) );
  DFFRX1 \bArray_reg[4][41]  ( .D(n6292), .CK(clk), .RN(n7587), .Q(
        \bArray[4][41] ), .QN(n5487) );
  DFFRX1 \bArray_reg[4][40]  ( .D(n6291), .CK(clk), .RN(n7587), .Q(
        \bArray[4][40] ), .QN(n5486) );
  DFFRX1 \bArray_reg[8][43]  ( .D(n6102), .CK(clk), .RN(n7603), .Q(
        \bArray[8][43] ), .QN(n5297) );
  DFFRX1 \bArray_reg[8][42]  ( .D(n6101), .CK(clk), .RN(n7603), .Q(
        \bArray[8][42] ), .QN(n5296) );
  DFFRX1 \bArray_reg[8][41]  ( .D(n6100), .CK(clk), .RN(n7603), .Q(
        \bArray[8][41] ), .QN(n5295) );
  DFFRX1 \bArray_reg[8][40]  ( .D(n6099), .CK(clk), .RN(n7603), .Q(
        \bArray[8][40] ), .QN(n5294) );
  DFFRX1 \bArray_reg[12][43]  ( .D(n5910), .CK(clk), .RN(n7619), .Q(
        \bArray[12][43] ), .QN(n5105) );
  DFFRX1 \bArray_reg[12][42]  ( .D(n5909), .CK(clk), .RN(n7619), .Q(
        \bArray[12][42] ), .QN(n5104) );
  DFFRX1 \bArray_reg[12][41]  ( .D(n5908), .CK(clk), .RN(n7619), .Q(
        \bArray[12][41] ), .QN(n5103) );
  DFFRX1 \bArray_reg[12][40]  ( .D(n5907), .CK(clk), .RN(n7619), .Q(
        \bArray[12][40] ), .QN(n5102) );
  DFFRX1 \bArray_reg[2][43]  ( .D(n6390), .CK(clk), .RN(n7579), .Q(
        \bArray[2][43] ), .QN(n5585) );
  DFFRX1 \bArray_reg[2][42]  ( .D(n6389), .CK(clk), .RN(n7579), .Q(
        \bArray[2][42] ), .QN(n5584) );
  DFFRX1 \bArray_reg[2][41]  ( .D(n6388), .CK(clk), .RN(n7579), .Q(
        \bArray[2][41] ), .QN(n5583) );
  DFFRX1 \bArray_reg[2][40]  ( .D(n6387), .CK(clk), .RN(n7579), .Q(
        \bArray[2][40] ), .QN(n5582) );
  DFFRX1 \bArray_reg[6][43]  ( .D(n6198), .CK(clk), .RN(n7595), .Q(
        \bArray[6][43] ), .QN(n5393) );
  DFFRX1 \bArray_reg[6][42]  ( .D(n6197), .CK(clk), .RN(n7595), .Q(
        \bArray[6][42] ), .QN(n5392) );
  DFFRX1 \bArray_reg[6][41]  ( .D(n6196), .CK(clk), .RN(n7595), .Q(
        \bArray[6][41] ), .QN(n5391) );
  DFFRX1 \bArray_reg[6][40]  ( .D(n6195), .CK(clk), .RN(n7595), .Q(
        \bArray[6][40] ), .QN(n5390) );
  DFFRX1 \bArray_reg[10][43]  ( .D(n6006), .CK(clk), .RN(n7611), .Q(
        \bArray[10][43] ), .QN(n5201) );
  DFFRX1 \bArray_reg[10][42]  ( .D(n6005), .CK(clk), .RN(n7611), .Q(
        \bArray[10][42] ), .QN(n5200) );
  DFFRX1 \bArray_reg[10][41]  ( .D(n6004), .CK(clk), .RN(n7611), .Q(
        \bArray[10][41] ), .QN(n5199) );
  DFFRX1 \bArray_reg[10][40]  ( .D(n6003), .CK(clk), .RN(n7611), .Q(
        \bArray[10][40] ), .QN(n5198) );
  DFFRX1 \bArray_reg[14][43]  ( .D(n5814), .CK(clk), .RN(n7627), .Q(
        \bArray[14][43] ), .QN(n5009) );
  DFFRX1 \bArray_reg[14][42]  ( .D(n5813), .CK(clk), .RN(n7627), .Q(
        \bArray[14][42] ), .QN(n5008) );
  DFFRX1 \bArray_reg[14][41]  ( .D(n5812), .CK(clk), .RN(n7627), .Q(
        \bArray[14][41] ), .QN(n5007) );
  DFFRX1 \bArray_reg[14][40]  ( .D(n5811), .CK(clk), .RN(n7627), .Q(
        \bArray[14][40] ), .QN(n5006) );
  DFFQX1 \xArray_reg[3][46]  ( .D(N28623), .CK(clk), .Q(\xArray[3][46] ) );
  DFFQX1 \xArray_reg[3][45]  ( .D(N28622), .CK(clk), .Q(\xArray[3][45] ) );
  DFFQX1 \xArray_reg[15][47]  ( .D(N27856), .CK(clk), .Q(\xArray[15][47] ) );
  DFFQX1 \xArray_reg[15][46]  ( .D(N27855), .CK(clk), .Q(\xArray[15][46] ) );
  DFFQX1 \xArray_reg[15][45]  ( .D(N27854), .CK(clk), .Q(\xArray[15][45] ) );
  DFFQX1 \xArray_reg[0][47]  ( .D(N28816), .CK(clk), .Q(\xArray[0][47] ) );
  DFFQX1 \xArray_reg[0][46]  ( .D(N28815), .CK(clk), .Q(\xArray[0][46] ) );
  DFFQX1 \xArray_reg[0][45]  ( .D(N28814), .CK(clk), .Q(\xArray[0][45] ) );
  DFFQX1 \xArray_reg[4][47]  ( .D(N28560), .CK(clk), .Q(\xArray[4][47] ) );
  DFFQX1 \xArray_reg[5][47]  ( .D(N28496), .CK(clk), .Q(\xArray[5][47] ) );
  DFFQX1 \xArray_reg[4][46]  ( .D(N28559), .CK(clk), .Q(\xArray[4][46] ) );
  DFFQX1 \xArray_reg[5][46]  ( .D(N28495), .CK(clk), .Q(\xArray[5][46] ) );
  DFFQX1 \xArray_reg[4][45]  ( .D(N28558), .CK(clk), .Q(\xArray[4][45] ) );
  DFFQX1 \xArray_reg[5][45]  ( .D(N28494), .CK(clk), .Q(\xArray[5][45] ) );
  DFFQX1 \xArray_reg[5][44]  ( .D(N28493), .CK(clk), .Q(\xArray[5][44] ) );
  DFFQX1 \xArray_reg[14][47]  ( .D(N27920), .CK(clk), .Q(\xArray[14][47] ) );
  DFFQX1 \xArray_reg[14][46]  ( .D(N27919), .CK(clk), .Q(\xArray[14][46] ) );
  DFFQX1 \xArray_reg[14][45]  ( .D(N27918), .CK(clk), .Q(\xArray[14][45] ) );
  DFFQX1 \xArray_reg[11][47]  ( .D(N28112), .CK(clk), .Q(\xArray[11][47] ) );
  DFFQX1 \xArray_reg[12][47]  ( .D(N28048), .CK(clk), .Q(\xArray[12][47] ) );
  DFFQX1 \xArray_reg[11][46]  ( .D(N28111), .CK(clk), .Q(\xArray[11][46] ) );
  DFFQX1 \xArray_reg[12][46]  ( .D(N28047), .CK(clk), .Q(\xArray[12][46] ) );
  DFFQX1 \xArray_reg[11][45]  ( .D(N28110), .CK(clk), .Q(\xArray[11][45] ) );
  DFFQX1 \xArray_reg[12][45]  ( .D(N28046), .CK(clk), .Q(\xArray[12][45] ) );
  DFFQX1 \xArray_reg[7][46]  ( .D(N28367), .CK(clk), .Q(\xArray[7][46] ) );
  DFFQX1 \xArray_reg[7][45]  ( .D(N28366), .CK(clk), .Q(\xArray[7][45] ) );
  DFFQX1 \xArray_reg[1][47]  ( .D(N28752), .CK(clk), .Q(\xArray[1][47] ) );
  DFFQX1 \xArray_reg[1][46]  ( .D(N28751), .CK(clk), .Q(\xArray[1][46] ) );
  DFFQX1 \xArray_reg[1][45]  ( .D(N28750), .CK(clk), .Q(\xArray[1][45] ) );
  DFFQX1 \xArray_reg[13][47]  ( .D(N27984), .CK(clk), .Q(\xArray[13][47] ) );
  DFFQX1 \xArray_reg[13][46]  ( .D(N27983), .CK(clk), .Q(\xArray[13][46] ) );
  DFFQX1 \xArray_reg[13][45]  ( .D(N27982), .CK(clk), .Q(\xArray[13][45] ) );
  DFFQX1 \xArray_reg[9][47]  ( .D(N28240), .CK(clk), .Q(\xArray[9][47] ) );
  DFFQX1 \xArray_reg[9][46]  ( .D(N28239), .CK(clk), .Q(\xArray[9][46] ) );
  DFFQX1 \xArray_reg[9][45]  ( .D(N28238), .CK(clk), .Q(\xArray[9][45] ) );
  DFFQX1 \xArray_reg[8][47]  ( .D(N28304), .CK(clk), .Q(\xArray[8][47] ) );
  DFFQX1 \xArray_reg[8][46]  ( .D(N28303), .CK(clk), .Q(\xArray[8][46] ) );
  DFFQX1 \xArray_reg[8][45]  ( .D(N28302), .CK(clk), .Q(\xArray[8][45] ) );
  DFFQX1 \xArray_reg[10][46]  ( .D(N28175), .CK(clk), .Q(\xArray[10][46] ) );
  DFFQX1 \xArray_reg[10][45]  ( .D(N28174), .CK(clk), .Q(\xArray[10][45] ) );
  DFFQX1 \xArray_reg[6][46]  ( .D(N28431), .CK(clk), .Q(\xArray[6][46] ) );
  DFFQX1 \xArray_reg[6][45]  ( .D(N28430), .CK(clk), .Q(\xArray[6][45] ) );
  DFFQX1 \xArray_reg[3][44]  ( .D(N28621), .CK(clk), .Q(\xArray[3][44] ) );
  DFFQX1 \xArray_reg[3][43]  ( .D(N28620), .CK(clk), .Q(\xArray[3][43] ) );
  DFFQX1 \xArray_reg[15][44]  ( .D(N27853), .CK(clk), .Q(\xArray[15][44] ) );
  DFFQX1 \xArray_reg[15][43]  ( .D(N27852), .CK(clk), .Q(\xArray[15][43] ) );
  DFFQX1 \xArray_reg[0][44]  ( .D(N28813), .CK(clk), .Q(\xArray[0][44] ) );
  DFFQX1 \xArray_reg[4][44]  ( .D(N28557), .CK(clk), .Q(\xArray[4][44] ) );
  DFFQX1 \xArray_reg[5][43]  ( .D(N28492), .CK(clk), .Q(\xArray[5][43] ) );
  DFFQX1 \xArray_reg[14][44]  ( .D(N27917), .CK(clk), .Q(\xArray[14][44] ) );
  DFFQX1 \xArray_reg[14][43]  ( .D(N27916), .CK(clk), .Q(\xArray[14][43] ) );
  DFFQX1 \xArray_reg[11][44]  ( .D(N28109), .CK(clk), .Q(\xArray[11][44] ) );
  DFFQX1 \xArray_reg[12][44]  ( .D(N28045), .CK(clk), .Q(\xArray[12][44] ) );
  DFFQX1 \xArray_reg[11][43]  ( .D(N28108), .CK(clk), .Q(\xArray[11][43] ) );
  DFFQX1 \xArray_reg[7][44]  ( .D(N28365), .CK(clk), .Q(\xArray[7][44] ) );
  DFFQX1 \xArray_reg[7][43]  ( .D(N28364), .CK(clk), .Q(\xArray[7][43] ) );
  DFFQX1 \xArray_reg[1][44]  ( .D(N28749), .CK(clk), .Q(\xArray[1][44] ) );
  DFFQX1 \xArray_reg[13][44]  ( .D(N27981), .CK(clk), .Q(\xArray[13][44] ) );
  DFFQX1 \xArray_reg[9][44]  ( .D(N28237), .CK(clk), .Q(\xArray[9][44] ) );
  DFFQX1 \xArray_reg[9][43]  ( .D(N28236), .CK(clk), .Q(\xArray[9][43] ) );
  DFFQX1 \xArray_reg[8][44]  ( .D(N28301), .CK(clk), .Q(\xArray[8][44] ) );
  DFFQX1 \xArray_reg[10][44]  ( .D(N28173), .CK(clk), .Q(\xArray[10][44] ) );
  DFFQX1 \xArray_reg[10][43]  ( .D(N28172), .CK(clk), .Q(\xArray[10][43] ) );
  DFFQX1 \xArray_reg[6][44]  ( .D(N28429), .CK(clk), .Q(\xArray[6][44] ) );
  DFFQX1 \xArray_reg[6][43]  ( .D(N28428), .CK(clk), .Q(\xArray[6][43] ) );
  DFFRX1 \bArray_reg[1][39]  ( .D(n6434), .CK(clk), .RN(n7576), .Q(
        \bArray[1][39] ), .QN(n5629) );
  DFFRX1 \bArray_reg[1][38]  ( .D(n6433), .CK(clk), .RN(n7576), .Q(
        \bArray[1][38] ), .QN(n5628) );
  DFFRX1 \bArray_reg[1][37]  ( .D(n6432), .CK(clk), .RN(n7576), .Q(
        \bArray[1][37] ), .QN(n5627) );
  DFFRX1 \bArray_reg[1][36]  ( .D(n6431), .CK(clk), .RN(n7576), .Q(
        \bArray[1][36] ), .QN(n5626) );
  DFFRX1 \bArray_reg[5][39]  ( .D(n6242), .CK(clk), .RN(n7592), .Q(
        \bArray[5][39] ), .QN(n5437) );
  DFFRX1 \bArray_reg[5][38]  ( .D(n6241), .CK(clk), .RN(n7592), .Q(
        \bArray[5][38] ), .QN(n5436) );
  DFFRX1 \bArray_reg[5][37]  ( .D(n6240), .CK(clk), .RN(n7592), .Q(
        \bArray[5][37] ), .QN(n5435) );
  DFFRX1 \bArray_reg[5][36]  ( .D(n6239), .CK(clk), .RN(n7592), .Q(
        \bArray[5][36] ), .QN(n5434) );
  DFFRX1 \bArray_reg[9][39]  ( .D(n6050), .CK(clk), .RN(n7608), .Q(
        \bArray[9][39] ), .QN(n5245) );
  DFFRX1 \bArray_reg[9][38]  ( .D(n6049), .CK(clk), .RN(n7608), .Q(
        \bArray[9][38] ), .QN(n5244) );
  DFFRX1 \bArray_reg[9][37]  ( .D(n6048), .CK(clk), .RN(n7608), .Q(
        \bArray[9][37] ), .QN(n5243) );
  DFFRX1 \bArray_reg[9][36]  ( .D(n6047), .CK(clk), .RN(n7608), .Q(
        \bArray[9][36] ), .QN(n5242) );
  DFFRX1 \bArray_reg[13][39]  ( .D(n5858), .CK(clk), .RN(n7624), .Q(
        \bArray[13][39] ), .QN(n5053) );
  DFFRX1 \bArray_reg[13][38]  ( .D(n5857), .CK(clk), .RN(n7624), .Q(
        \bArray[13][38] ), .QN(n5052) );
  DFFRX1 \bArray_reg[13][37]  ( .D(n5856), .CK(clk), .RN(n7624), .Q(
        \bArray[13][37] ), .QN(n5051) );
  DFFRX1 \bArray_reg[13][36]  ( .D(n5855), .CK(clk), .RN(n7624), .Q(
        \bArray[13][36] ), .QN(n5050) );
  DFFRX1 \bArray_reg[3][39]  ( .D(n6338), .CK(clk), .RN(n7584), .Q(
        \bArray[3][39] ), .QN(n5533) );
  DFFRX1 \bArray_reg[3][38]  ( .D(n6337), .CK(clk), .RN(n7584), .Q(
        \bArray[3][38] ), .QN(n5532) );
  DFFRX1 \bArray_reg[3][37]  ( .D(n6336), .CK(clk), .RN(n7584), .Q(
        \bArray[3][37] ), .QN(n5531) );
  DFFRX1 \bArray_reg[3][36]  ( .D(n6335), .CK(clk), .RN(n7584), .Q(
        \bArray[3][36] ), .QN(n5530) );
  DFFRX1 \bArray_reg[7][39]  ( .D(n6146), .CK(clk), .RN(n7600), .Q(
        \bArray[7][39] ), .QN(n5341) );
  DFFRX1 \bArray_reg[7][38]  ( .D(n6145), .CK(clk), .RN(n7600), .Q(
        \bArray[7][38] ), .QN(n5340) );
  DFFRX1 \bArray_reg[7][37]  ( .D(n6144), .CK(clk), .RN(n7600), .Q(
        \bArray[7][37] ), .QN(n5339) );
  DFFRX1 \bArray_reg[7][36]  ( .D(n6143), .CK(clk), .RN(n7600), .Q(
        \bArray[7][36] ), .QN(n5338) );
  DFFRX1 \bArray_reg[11][39]  ( .D(n5954), .CK(clk), .RN(n7616), .Q(
        \bArray[11][39] ), .QN(n5149) );
  DFFRX1 \bArray_reg[11][38]  ( .D(n5953), .CK(clk), .RN(n7616), .Q(
        \bArray[11][38] ), .QN(n5148) );
  DFFRX1 \bArray_reg[11][37]  ( .D(n5952), .CK(clk), .RN(n7616), .Q(
        \bArray[11][37] ), .QN(n5147) );
  DFFRX1 \bArray_reg[11][36]  ( .D(n5951), .CK(clk), .RN(n7616), .Q(
        \bArray[11][36] ), .QN(n5146) );
  DFFRX1 \bArray_reg[15][39]  ( .D(n5762), .CK(clk), .RN(n7632), .Q(
        \bArray[15][39] ), .QN(n4957) );
  DFFRX1 \bArray_reg[15][38]  ( .D(n5761), .CK(clk), .RN(n7632), .Q(
        \bArray[15][38] ), .QN(n4956) );
  DFFRX1 \bArray_reg[15][37]  ( .D(n5760), .CK(clk), .RN(n7632), .Q(
        \bArray[15][37] ), .QN(n4955) );
  DFFRX1 \bArray_reg[15][36]  ( .D(n5759), .CK(clk), .RN(n7632), .Q(
        \bArray[15][36] ), .QN(n4954) );
  DFFRX1 \bArray_reg[0][39]  ( .D(n6482), .CK(clk), .RN(n7572), .Q(
        \bArray[0][39] ), .QN(n5677) );
  DFFRX1 \bArray_reg[0][38]  ( .D(n6481), .CK(clk), .RN(n7572), .Q(
        \bArray[0][38] ), .QN(n5676) );
  DFFRX1 \bArray_reg[0][37]  ( .D(n6480), .CK(clk), .RN(n7572), .Q(
        \bArray[0][37] ), .QN(n5675) );
  DFFRX1 \bArray_reg[0][36]  ( .D(n6479), .CK(clk), .RN(n7572), .Q(
        \bArray[0][36] ), .QN(n5674) );
  DFFRX1 \bArray_reg[4][39]  ( .D(n6290), .CK(clk), .RN(n7588), .Q(
        \bArray[4][39] ), .QN(n5485) );
  DFFRX1 \bArray_reg[4][38]  ( .D(n6289), .CK(clk), .RN(n7588), .Q(
        \bArray[4][38] ), .QN(n5484) );
  DFFRX1 \bArray_reg[4][37]  ( .D(n6288), .CK(clk), .RN(n7588), .Q(
        \bArray[4][37] ), .QN(n5483) );
  DFFRX1 \bArray_reg[4][36]  ( .D(n6287), .CK(clk), .RN(n7588), .Q(
        \bArray[4][36] ), .QN(n5482) );
  DFFRX1 \bArray_reg[8][39]  ( .D(n6098), .CK(clk), .RN(n7604), .Q(
        \bArray[8][39] ), .QN(n5293) );
  DFFRX1 \bArray_reg[8][38]  ( .D(n6097), .CK(clk), .RN(n7604), .Q(
        \bArray[8][38] ), .QN(n5292) );
  DFFRX1 \bArray_reg[8][37]  ( .D(n6096), .CK(clk), .RN(n7604), .Q(
        \bArray[8][37] ), .QN(n5291) );
  DFFRX1 \bArray_reg[8][36]  ( .D(n6095), .CK(clk), .RN(n7604), .Q(
        \bArray[8][36] ), .QN(n5290) );
  DFFRX1 \bArray_reg[12][39]  ( .D(n5906), .CK(clk), .RN(n7620), .Q(
        \bArray[12][39] ), .QN(n5101) );
  DFFRX1 \bArray_reg[12][38]  ( .D(n5905), .CK(clk), .RN(n7620), .Q(
        \bArray[12][38] ), .QN(n5100) );
  DFFRX1 \bArray_reg[12][37]  ( .D(n5904), .CK(clk), .RN(n7620), .Q(
        \bArray[12][37] ), .QN(n5099) );
  DFFRX1 \bArray_reg[12][36]  ( .D(n5903), .CK(clk), .RN(n7620), .Q(
        \bArray[12][36] ), .QN(n5098) );
  DFFRX1 \bArray_reg[2][39]  ( .D(n6386), .CK(clk), .RN(n7580), .Q(
        \bArray[2][39] ), .QN(n5581) );
  DFFRX1 \bArray_reg[2][38]  ( .D(n6385), .CK(clk), .RN(n7580), .Q(
        \bArray[2][38] ), .QN(n5580) );
  DFFRX1 \bArray_reg[2][37]  ( .D(n6384), .CK(clk), .RN(n7580), .Q(
        \bArray[2][37] ), .QN(n5579) );
  DFFRX1 \bArray_reg[2][36]  ( .D(n6383), .CK(clk), .RN(n7580), .Q(
        \bArray[2][36] ), .QN(n5578) );
  DFFRX1 \bArray_reg[6][39]  ( .D(n6194), .CK(clk), .RN(n7596), .Q(
        \bArray[6][39] ), .QN(n5389) );
  DFFRX1 \bArray_reg[6][38]  ( .D(n6193), .CK(clk), .RN(n7596), .Q(
        \bArray[6][38] ), .QN(n5388) );
  DFFRX1 \bArray_reg[6][37]  ( .D(n6192), .CK(clk), .RN(n7596), .Q(
        \bArray[6][37] ), .QN(n5387) );
  DFFRX1 \bArray_reg[6][36]  ( .D(n6191), .CK(clk), .RN(n7596), .Q(
        \bArray[6][36] ), .QN(n5386) );
  DFFRX1 \bArray_reg[10][39]  ( .D(n6002), .CK(clk), .RN(n7612), .Q(
        \bArray[10][39] ), .QN(n5197) );
  DFFRX1 \bArray_reg[10][38]  ( .D(n6001), .CK(clk), .RN(n7612), .Q(
        \bArray[10][38] ), .QN(n5196) );
  DFFRX1 \bArray_reg[10][37]  ( .D(n6000), .CK(clk), .RN(n7612), .Q(
        \bArray[10][37] ), .QN(n5195) );
  DFFRX1 \bArray_reg[10][36]  ( .D(n5999), .CK(clk), .RN(n7612), .Q(
        \bArray[10][36] ), .QN(n5194) );
  DFFRX1 \bArray_reg[14][39]  ( .D(n5810), .CK(clk), .RN(n7628), .Q(
        \bArray[14][39] ), .QN(n5005) );
  DFFRX1 \bArray_reg[14][38]  ( .D(n5809), .CK(clk), .RN(n7628), .Q(
        \bArray[14][38] ), .QN(n5004) );
  DFFRX1 \bArray_reg[14][37]  ( .D(n5808), .CK(clk), .RN(n7628), .Q(
        \bArray[14][37] ), .QN(n5003) );
  DFFRX1 \bArray_reg[14][36]  ( .D(n5807), .CK(clk), .RN(n7628), .Q(
        \bArray[14][36] ), .QN(n5002) );
  DFFQX1 \xArray_reg[3][42]  ( .D(N28619), .CK(clk), .Q(\xArray[3][42] ) );
  DFFQX1 \xArray_reg[15][42]  ( .D(N27851), .CK(clk), .Q(\xArray[15][42] ) );
  DFFQX1 \xArray_reg[0][43]  ( .D(N28812), .CK(clk), .Q(\xArray[0][43] ) );
  DFFQX1 \xArray_reg[0][42]  ( .D(N28811), .CK(clk), .Q(\xArray[0][42] ) );
  DFFQX1 \xArray_reg[4][43]  ( .D(N28556), .CK(clk), .Q(\xArray[4][43] ) );
  DFFQX1 \xArray_reg[4][42]  ( .D(N28555), .CK(clk), .Q(\xArray[4][42] ) );
  DFFQX1 \xArray_reg[5][42]  ( .D(N28491), .CK(clk), .Q(\xArray[5][42] ) );
  DFFQX1 \xArray_reg[14][42]  ( .D(N27915), .CK(clk), .Q(\xArray[14][42] ) );
  DFFQX1 \xArray_reg[12][43]  ( .D(N28044), .CK(clk), .Q(\xArray[12][43] ) );
  DFFQX1 \xArray_reg[11][42]  ( .D(N28107), .CK(clk), .Q(\xArray[11][42] ) );
  DFFQX1 \xArray_reg[12][42]  ( .D(N28043), .CK(clk), .Q(\xArray[12][42] ) );
  DFFQX1 \xArray_reg[7][42]  ( .D(N28363), .CK(clk), .Q(\xArray[7][42] ) );
  DFFQX1 \xArray_reg[1][43]  ( .D(N28748), .CK(clk), .Q(\xArray[1][43] ) );
  DFFQX1 \xArray_reg[1][42]  ( .D(N28747), .CK(clk), .Q(\xArray[1][42] ) );
  DFFQX1 \xArray_reg[13][43]  ( .D(N27980), .CK(clk), .Q(\xArray[13][43] ) );
  DFFQX1 \xArray_reg[13][42]  ( .D(N27979), .CK(clk), .Q(\xArray[13][42] ) );
  DFFQX1 \xArray_reg[9][42]  ( .D(N28235), .CK(clk), .Q(\xArray[9][42] ) );
  DFFQX1 \xArray_reg[8][43]  ( .D(N28300), .CK(clk), .Q(\xArray[8][43] ) );
  DFFQX1 \xArray_reg[8][42]  ( .D(N28299), .CK(clk), .Q(\xArray[8][42] ) );
  DFFQX1 \xArray_reg[10][42]  ( .D(N28171), .CK(clk), .Q(\xArray[10][42] ) );
  DFFQX1 \xArray_reg[10][41]  ( .D(N28170), .CK(clk), .Q(\xArray[10][41] ) );
  DFFQX1 \xArray_reg[6][42]  ( .D(N28427), .CK(clk), .Q(\xArray[6][42] ) );
  DFFQX1 \xArray_reg[6][41]  ( .D(N28426), .CK(clk), .Q(\xArray[6][41] ) );
  DFFQX1 \xArray_reg[1][41]  ( .D(N28746), .CK(clk), .Q(\xArray[1][41] ) );
  DFFQX1 \xArray_reg[1][40]  ( .D(N28745), .CK(clk), .Q(\xArray[1][40] ) );
  DFFQX1 \xArray_reg[13][41]  ( .D(N27978), .CK(clk), .Q(\xArray[13][41] ) );
  DFFQX1 \xArray_reg[13][40]  ( .D(N27977), .CK(clk), .Q(\xArray[13][40] ) );
  DFFQX1 \xArray_reg[9][41]  ( .D(N28234), .CK(clk), .Q(\xArray[9][41] ) );
  DFFQX1 \xArray_reg[9][40]  ( .D(N28233), .CK(clk), .Q(\xArray[9][40] ) );
  DFFQX1 \xArray_reg[8][41]  ( .D(N28298), .CK(clk), .Q(\xArray[8][41] ) );
  DFFQX1 \xArray_reg[8][40]  ( .D(N28297), .CK(clk), .Q(\xArray[8][40] ) );
  DFFQX1 \xArray_reg[10][40]  ( .D(N28169), .CK(clk), .Q(\xArray[10][40] ) );
  DFFQX1 \xArray_reg[10][39]  ( .D(N28168), .CK(clk), .Q(\xArray[10][39] ) );
  DFFQX1 \xArray_reg[6][40]  ( .D(N28425), .CK(clk), .Q(\xArray[6][40] ) );
  DFFQX1 \xArray_reg[6][39]  ( .D(N28424), .CK(clk), .Q(\xArray[6][39] ) );
  DFFRX1 \bArray_reg[1][35]  ( .D(n6430), .CK(clk), .RN(n7576), .Q(
        \bArray[1][35] ), .QN(n5625) );
  DFFRX1 \bArray_reg[1][34]  ( .D(n6429), .CK(clk), .RN(n7576), .Q(
        \bArray[1][34] ), .QN(n5624) );
  DFFRX1 \bArray_reg[1][33]  ( .D(n6428), .CK(clk), .RN(n7576), .Q(
        \bArray[1][33] ), .QN(n5623) );
  DFFRX1 \bArray_reg[1][32]  ( .D(n6427), .CK(clk), .RN(n7576), .Q(
        \bArray[1][32] ), .QN(n5622) );
  DFFRX1 \bArray_reg[5][35]  ( .D(n6238), .CK(clk), .RN(n7592), .Q(
        \bArray[5][35] ), .QN(n5433) );
  DFFRX1 \bArray_reg[5][34]  ( .D(n6237), .CK(clk), .RN(n7592), .Q(
        \bArray[5][34] ), .QN(n5432) );
  DFFRX1 \bArray_reg[5][33]  ( .D(n6236), .CK(clk), .RN(n7592), .Q(
        \bArray[5][33] ), .QN(n5431) );
  DFFRX1 \bArray_reg[5][32]  ( .D(n6235), .CK(clk), .RN(n7592), .Q(
        \bArray[5][32] ), .QN(n5430) );
  DFFRX1 \bArray_reg[9][35]  ( .D(n6046), .CK(clk), .RN(n7608), .Q(
        \bArray[9][35] ), .QN(n5241) );
  DFFRX1 \bArray_reg[9][34]  ( .D(n6045), .CK(clk), .RN(n7608), .Q(
        \bArray[9][34] ), .QN(n5240) );
  DFFRX1 \bArray_reg[9][33]  ( .D(n6044), .CK(clk), .RN(n7608), .Q(
        \bArray[9][33] ), .QN(n5239) );
  DFFRX1 \bArray_reg[9][32]  ( .D(n6043), .CK(clk), .RN(n7608), .Q(
        \bArray[9][32] ), .QN(n5238) );
  DFFRX1 \bArray_reg[13][35]  ( .D(n5854), .CK(clk), .RN(n7624), .Q(
        \bArray[13][35] ), .QN(n5049) );
  DFFRX1 \bArray_reg[13][34]  ( .D(n5853), .CK(clk), .RN(n7624), .Q(
        \bArray[13][34] ), .QN(n5048) );
  DFFRX1 \bArray_reg[13][33]  ( .D(n5852), .CK(clk), .RN(n7624), .Q(
        \bArray[13][33] ), .QN(n5047) );
  DFFRX1 \bArray_reg[13][32]  ( .D(n5851), .CK(clk), .RN(n7624), .Q(
        \bArray[13][32] ), .QN(n5046) );
  DFFRX1 \bArray_reg[3][35]  ( .D(n6334), .CK(clk), .RN(n7584), .Q(
        \bArray[3][35] ), .QN(n5529) );
  DFFRX1 \bArray_reg[3][34]  ( .D(n6333), .CK(clk), .RN(n7584), .Q(
        \bArray[3][34] ), .QN(n5528) );
  DFFRX1 \bArray_reg[3][33]  ( .D(n6332), .CK(clk), .RN(n7584), .Q(
        \bArray[3][33] ), .QN(n5527) );
  DFFRX1 \bArray_reg[3][32]  ( .D(n6331), .CK(clk), .RN(n7584), .Q(
        \bArray[3][32] ), .QN(n5526) );
  DFFRX1 \bArray_reg[7][35]  ( .D(n6142), .CK(clk), .RN(n7600), .Q(
        \bArray[7][35] ), .QN(n5337) );
  DFFRX1 \bArray_reg[7][34]  ( .D(n6141), .CK(clk), .RN(n7600), .Q(
        \bArray[7][34] ), .QN(n5336) );
  DFFRX1 \bArray_reg[7][33]  ( .D(n6140), .CK(clk), .RN(n7600), .Q(
        \bArray[7][33] ), .QN(n5335) );
  DFFRX1 \bArray_reg[7][32]  ( .D(n6139), .CK(clk), .RN(n7600), .Q(
        \bArray[7][32] ), .QN(n5334) );
  DFFRX1 \bArray_reg[11][35]  ( .D(n5950), .CK(clk), .RN(n7616), .Q(
        \bArray[11][35] ), .QN(n5145) );
  DFFRX1 \bArray_reg[11][34]  ( .D(n5949), .CK(clk), .RN(n7616), .Q(
        \bArray[11][34] ), .QN(n5144) );
  DFFRX1 \bArray_reg[11][33]  ( .D(n5948), .CK(clk), .RN(n7616), .Q(
        \bArray[11][33] ), .QN(n5143) );
  DFFRX1 \bArray_reg[11][32]  ( .D(n5947), .CK(clk), .RN(n7616), .Q(
        \bArray[11][32] ), .QN(n5142) );
  DFFRX1 \bArray_reg[15][35]  ( .D(n5758), .CK(clk), .RN(n7632), .Q(
        \bArray[15][35] ), .QN(n4953) );
  DFFRX1 \bArray_reg[15][34]  ( .D(n5757), .CK(clk), .RN(n7632), .Q(
        \bArray[15][34] ), .QN(n4952) );
  DFFRX1 \bArray_reg[15][33]  ( .D(n5756), .CK(clk), .RN(n7632), .Q(
        \bArray[15][33] ), .QN(n4951) );
  DFFRX1 \bArray_reg[15][32]  ( .D(n5755), .CK(clk), .RN(n7632), .Q(
        \bArray[15][32] ), .QN(n4950) );
  DFFRX1 \bArray_reg[0][35]  ( .D(n6478), .CK(clk), .RN(n7572), .Q(
        \bArray[0][35] ), .QN(n5673) );
  DFFRX1 \bArray_reg[0][34]  ( .D(n6477), .CK(clk), .RN(n7572), .Q(
        \bArray[0][34] ), .QN(n5672) );
  DFFRX1 \bArray_reg[0][33]  ( .D(n6476), .CK(clk), .RN(n7572), .Q(
        \bArray[0][33] ), .QN(n5671) );
  DFFRX1 \bArray_reg[0][32]  ( .D(n6475), .CK(clk), .RN(n7572), .Q(
        \bArray[0][32] ), .QN(n5670) );
  DFFRX1 \bArray_reg[4][35]  ( .D(n6286), .CK(clk), .RN(n7588), .Q(
        \bArray[4][35] ), .QN(n5481) );
  DFFRX1 \bArray_reg[4][34]  ( .D(n6285), .CK(clk), .RN(n7588), .Q(
        \bArray[4][34] ), .QN(n5480) );
  DFFRX1 \bArray_reg[4][33]  ( .D(n6284), .CK(clk), .RN(n7588), .Q(
        \bArray[4][33] ), .QN(n5479) );
  DFFRX1 \bArray_reg[4][32]  ( .D(n6283), .CK(clk), .RN(n7588), .Q(
        \bArray[4][32] ), .QN(n5478) );
  DFFRX1 \bArray_reg[8][35]  ( .D(n6094), .CK(clk), .RN(n7604), .Q(
        \bArray[8][35] ), .QN(n5289) );
  DFFRX1 \bArray_reg[8][34]  ( .D(n6093), .CK(clk), .RN(n7604), .Q(
        \bArray[8][34] ), .QN(n5288) );
  DFFRX1 \bArray_reg[8][33]  ( .D(n6092), .CK(clk), .RN(n7604), .Q(
        \bArray[8][33] ), .QN(n5287) );
  DFFRX1 \bArray_reg[8][32]  ( .D(n6091), .CK(clk), .RN(n7604), .Q(
        \bArray[8][32] ), .QN(n5286) );
  DFFRX1 \bArray_reg[12][35]  ( .D(n5902), .CK(clk), .RN(n7620), .Q(
        \bArray[12][35] ), .QN(n5097) );
  DFFRX1 \bArray_reg[12][34]  ( .D(n5901), .CK(clk), .RN(n7620), .Q(
        \bArray[12][34] ), .QN(n5096) );
  DFFRX1 \bArray_reg[12][33]  ( .D(n5900), .CK(clk), .RN(n7620), .Q(
        \bArray[12][33] ), .QN(n5095) );
  DFFRX1 \bArray_reg[12][32]  ( .D(n5899), .CK(clk), .RN(n7620), .Q(
        \bArray[12][32] ), .QN(n5094) );
  DFFRX1 \bArray_reg[2][35]  ( .D(n6382), .CK(clk), .RN(n7580), .Q(
        \bArray[2][35] ), .QN(n5577) );
  DFFRX1 \bArray_reg[2][34]  ( .D(n6381), .CK(clk), .RN(n7580), .Q(
        \bArray[2][34] ), .QN(n5576) );
  DFFRX1 \bArray_reg[2][33]  ( .D(n6380), .CK(clk), .RN(n7580), .Q(
        \bArray[2][33] ), .QN(n5575) );
  DFFRX1 \bArray_reg[2][32]  ( .D(n6379), .CK(clk), .RN(n7580), .Q(
        \bArray[2][32] ), .QN(n5574) );
  DFFRX1 \bArray_reg[6][35]  ( .D(n6190), .CK(clk), .RN(n7596), .Q(
        \bArray[6][35] ), .QN(n5385) );
  DFFRX1 \bArray_reg[6][34]  ( .D(n6189), .CK(clk), .RN(n7596), .Q(
        \bArray[6][34] ), .QN(n5384) );
  DFFRX1 \bArray_reg[6][33]  ( .D(n6188), .CK(clk), .RN(n7596), .Q(
        \bArray[6][33] ), .QN(n5383) );
  DFFRX1 \bArray_reg[6][32]  ( .D(n6187), .CK(clk), .RN(n7596), .Q(
        \bArray[6][32] ), .QN(n5382) );
  DFFRX1 \bArray_reg[10][35]  ( .D(n5998), .CK(clk), .RN(n7612), .Q(
        \bArray[10][35] ), .QN(n5193) );
  DFFRX1 \bArray_reg[10][34]  ( .D(n5997), .CK(clk), .RN(n7612), .Q(
        \bArray[10][34] ), .QN(n5192) );
  DFFRX1 \bArray_reg[10][33]  ( .D(n5996), .CK(clk), .RN(n7612), .Q(
        \bArray[10][33] ), .QN(n5191) );
  DFFRX1 \bArray_reg[10][32]  ( .D(n5995), .CK(clk), .RN(n7612), .Q(
        \bArray[10][32] ), .QN(n5190) );
  DFFRX1 \bArray_reg[14][35]  ( .D(n5806), .CK(clk), .RN(n7628), .Q(
        \bArray[14][35] ), .QN(n5001) );
  DFFRX1 \bArray_reg[14][34]  ( .D(n5805), .CK(clk), .RN(n7628), .Q(
        \bArray[14][34] ), .QN(n5000) );
  DFFRX1 \bArray_reg[14][33]  ( .D(n5804), .CK(clk), .RN(n7628), .Q(
        \bArray[14][33] ), .QN(n4999) );
  DFFRX1 \bArray_reg[14][32]  ( .D(n5803), .CK(clk), .RN(n7628), .Q(
        \bArray[14][32] ), .QN(n4998) );
  DFFQX1 \xArray_reg[1][39]  ( .D(N28744), .CK(clk), .Q(\xArray[1][39] ) );
  DFFQX1 \xArray_reg[1][38]  ( .D(N28743), .CK(clk), .Q(\xArray[1][38] ) );
  DFFQX1 \xArray_reg[13][39]  ( .D(N27976), .CK(clk), .Q(\xArray[13][39] ) );
  DFFQX1 \xArray_reg[13][38]  ( .D(N27975), .CK(clk), .Q(\xArray[13][38] ) );
  DFFQX1 \xArray_reg[9][39]  ( .D(N28232), .CK(clk), .Q(\xArray[9][39] ) );
  DFFQX1 \xArray_reg[9][38]  ( .D(N28231), .CK(clk), .Q(\xArray[9][38] ) );
  DFFQX1 \xArray_reg[8][39]  ( .D(N28296), .CK(clk), .Q(\xArray[8][39] ) );
  DFFQX1 \xArray_reg[8][38]  ( .D(N28295), .CK(clk), .Q(\xArray[8][38] ) );
  DFFQX1 \xArray_reg[10][38]  ( .D(N28167), .CK(clk), .Q(\xArray[10][38] ) );
  DFFQX1 \xArray_reg[10][37]  ( .D(N28166), .CK(clk), .Q(\xArray[10][37] ) );
  DFFQX1 \xArray_reg[6][38]  ( .D(N28423), .CK(clk), .Q(\xArray[6][38] ) );
  DFFQX1 \xArray_reg[6][37]  ( .D(N28422), .CK(clk), .Q(\xArray[6][37] ) );
  DFFQX1 \xArray_reg[1][37]  ( .D(N28742), .CK(clk), .Q(\xArray[1][37] ) );
  DFFQX1 \xArray_reg[1][36]  ( .D(N28741), .CK(clk), .Q(\xArray[1][36] ) );
  DFFQX1 \xArray_reg[1][35]  ( .D(N28740), .CK(clk), .Q(\xArray[1][35] ) );
  DFFQX1 \xArray_reg[13][37]  ( .D(N27974), .CK(clk), .Q(\xArray[13][37] ) );
  DFFQX1 \xArray_reg[13][36]  ( .D(N27973), .CK(clk), .Q(\xArray[13][36] ) );
  DFFQX1 \xArray_reg[13][35]  ( .D(N27972), .CK(clk), .Q(\xArray[13][35] ) );
  DFFQX1 \xArray_reg[9][37]  ( .D(N28230), .CK(clk), .Q(\xArray[9][37] ) );
  DFFQX1 \xArray_reg[9][36]  ( .D(N28229), .CK(clk), .Q(\xArray[9][36] ) );
  DFFQX1 \xArray_reg[9][35]  ( .D(N28228), .CK(clk), .Q(\xArray[9][35] ) );
  DFFQX1 \xArray_reg[8][37]  ( .D(N28294), .CK(clk), .Q(\xArray[8][37] ) );
  DFFQX1 \xArray_reg[8][36]  ( .D(N28293), .CK(clk), .Q(\xArray[8][36] ) );
  DFFQX1 \xArray_reg[8][35]  ( .D(N28292), .CK(clk), .Q(\xArray[8][35] ) );
  DFFQX1 \xArray_reg[10][36]  ( .D(N28165), .CK(clk), .Q(\xArray[10][36] ) );
  DFFQX1 \xArray_reg[10][35]  ( .D(N28164), .CK(clk), .Q(\xArray[10][35] ) );
  DFFQX1 \xArray_reg[6][36]  ( .D(N28421), .CK(clk), .Q(\xArray[6][36] ) );
  DFFQX1 \xArray_reg[6][35]  ( .D(N28420), .CK(clk), .Q(\xArray[6][35] ) );
  DFFRX1 \bArray_reg[1][31]  ( .D(n6426), .CK(clk), .RN(n7576), .Q(
        \bArray[1][31] ), .QN(n5621) );
  DFFRX1 \bArray_reg[1][30]  ( .D(n6425), .CK(clk), .RN(n7576), .Q(
        \bArray[1][30] ), .QN(n5620) );
  DFFRX1 \bArray_reg[1][29]  ( .D(n6424), .CK(clk), .RN(n7576), .Q(
        \bArray[1][29] ), .QN(n5619) );
  DFFRX1 \bArray_reg[1][28]  ( .D(n6423), .CK(clk), .RN(n7576), .Q(
        \bArray[1][28] ), .QN(n5618) );
  DFFRX1 \bArray_reg[5][31]  ( .D(n6234), .CK(clk), .RN(n7592), .Q(
        \bArray[5][31] ), .QN(n5429) );
  DFFRX1 \bArray_reg[5][30]  ( .D(n6233), .CK(clk), .RN(n7592), .Q(
        \bArray[5][30] ), .QN(n5428) );
  DFFRX1 \bArray_reg[5][29]  ( .D(n6232), .CK(clk), .RN(n7592), .Q(
        \bArray[5][29] ), .QN(n5427) );
  DFFRX1 \bArray_reg[5][28]  ( .D(n6231), .CK(clk), .RN(n7592), .Q(
        \bArray[5][28] ), .QN(n5426) );
  DFFRX1 \bArray_reg[9][31]  ( .D(n6042), .CK(clk), .RN(n7608), .Q(
        \bArray[9][31] ), .QN(n5237) );
  DFFRX1 \bArray_reg[9][30]  ( .D(n6041), .CK(clk), .RN(n7608), .Q(
        \bArray[9][30] ), .QN(n5236) );
  DFFRX1 \bArray_reg[9][29]  ( .D(n6040), .CK(clk), .RN(n7608), .Q(
        \bArray[9][29] ), .QN(n5235) );
  DFFRX1 \bArray_reg[9][28]  ( .D(n6039), .CK(clk), .RN(n7608), .Q(
        \bArray[9][28] ), .QN(n5234) );
  DFFRX1 \bArray_reg[13][31]  ( .D(n5850), .CK(clk), .RN(n7624), .Q(
        \bArray[13][31] ), .QN(n5045) );
  DFFRX1 \bArray_reg[13][30]  ( .D(n5849), .CK(clk), .RN(n7624), .Q(
        \bArray[13][30] ), .QN(n5044) );
  DFFRX1 \bArray_reg[13][29]  ( .D(n5848), .CK(clk), .RN(n7624), .Q(
        \bArray[13][29] ), .QN(n5043) );
  DFFRX1 \bArray_reg[13][28]  ( .D(n5847), .CK(clk), .RN(n7624), .Q(
        \bArray[13][28] ), .QN(n5042) );
  DFFRX1 \bArray_reg[3][31]  ( .D(n6330), .CK(clk), .RN(n7584), .Q(
        \bArray[3][31] ), .QN(n5525) );
  DFFRX1 \bArray_reg[3][30]  ( .D(n6329), .CK(clk), .RN(n7584), .Q(
        \bArray[3][30] ), .QN(n5524) );
  DFFRX1 \bArray_reg[3][29]  ( .D(n6328), .CK(clk), .RN(n7584), .Q(
        \bArray[3][29] ), .QN(n5523) );
  DFFRX1 \bArray_reg[3][28]  ( .D(n6327), .CK(clk), .RN(n7584), .Q(
        \bArray[3][28] ), .QN(n5522) );
  DFFRX1 \bArray_reg[7][31]  ( .D(n6138), .CK(clk), .RN(n7600), .Q(
        \bArray[7][31] ), .QN(n5333) );
  DFFRX1 \bArray_reg[7][30]  ( .D(n6137), .CK(clk), .RN(n7600), .Q(
        \bArray[7][30] ), .QN(n5332) );
  DFFRX1 \bArray_reg[7][29]  ( .D(n6136), .CK(clk), .RN(n7600), .Q(
        \bArray[7][29] ), .QN(n5331) );
  DFFRX1 \bArray_reg[7][28]  ( .D(n6135), .CK(clk), .RN(n7600), .Q(
        \bArray[7][28] ), .QN(n5330) );
  DFFRX1 \bArray_reg[11][31]  ( .D(n5946), .CK(clk), .RN(n7616), .Q(
        \bArray[11][31] ), .QN(n5141) );
  DFFRX1 \bArray_reg[11][30]  ( .D(n5945), .CK(clk), .RN(n7616), .Q(
        \bArray[11][30] ), .QN(n5140) );
  DFFRX1 \bArray_reg[11][29]  ( .D(n5944), .CK(clk), .RN(n7616), .Q(
        \bArray[11][29] ), .QN(n5139) );
  DFFRX1 \bArray_reg[11][28]  ( .D(n5943), .CK(clk), .RN(n7616), .Q(
        \bArray[11][28] ), .QN(n5138) );
  DFFRX1 \bArray_reg[15][31]  ( .D(n5754), .CK(clk), .RN(n7632), .Q(
        \bArray[15][31] ), .QN(n4949) );
  DFFRX1 \bArray_reg[15][30]  ( .D(n5753), .CK(clk), .RN(n7632), .Q(
        \bArray[15][30] ), .QN(n4948) );
  DFFRX1 \bArray_reg[15][29]  ( .D(n5752), .CK(clk), .RN(n7632), .Q(
        \bArray[15][29] ), .QN(n4947) );
  DFFRX1 \bArray_reg[15][28]  ( .D(n5751), .CK(clk), .RN(n7632), .Q(
        \bArray[15][28] ), .QN(n4946) );
  DFFRX1 \bArray_reg[0][31]  ( .D(n6474), .CK(clk), .RN(n7572), .Q(
        \bArray[0][31] ), .QN(n5669) );
  DFFRX1 \bArray_reg[0][30]  ( .D(n6473), .CK(clk), .RN(n7572), .Q(
        \bArray[0][30] ), .QN(n5668) );
  DFFRX1 \bArray_reg[0][29]  ( .D(n6472), .CK(clk), .RN(n7572), .Q(
        \bArray[0][29] ), .QN(n5667) );
  DFFRX1 \bArray_reg[0][28]  ( .D(n6471), .CK(clk), .RN(n7572), .Q(
        \bArray[0][28] ), .QN(n5666) );
  DFFRX1 \bArray_reg[4][31]  ( .D(n6282), .CK(clk), .RN(n7588), .Q(
        \bArray[4][31] ), .QN(n5477) );
  DFFRX1 \bArray_reg[4][30]  ( .D(n6281), .CK(clk), .RN(n7588), .Q(
        \bArray[4][30] ), .QN(n5476) );
  DFFRX1 \bArray_reg[4][29]  ( .D(n6280), .CK(clk), .RN(n7588), .Q(
        \bArray[4][29] ), .QN(n5475) );
  DFFRX1 \bArray_reg[4][28]  ( .D(n6279), .CK(clk), .RN(n7588), .Q(
        \bArray[4][28] ), .QN(n5474) );
  DFFRX1 \bArray_reg[8][31]  ( .D(n6090), .CK(clk), .RN(n7604), .Q(
        \bArray[8][31] ), .QN(n5285) );
  DFFRX1 \bArray_reg[8][30]  ( .D(n6089), .CK(clk), .RN(n7604), .Q(
        \bArray[8][30] ), .QN(n5284) );
  DFFRX1 \bArray_reg[8][29]  ( .D(n6088), .CK(clk), .RN(n7604), .Q(
        \bArray[8][29] ), .QN(n5283) );
  DFFRX1 \bArray_reg[8][28]  ( .D(n6087), .CK(clk), .RN(n7604), .Q(
        \bArray[8][28] ), .QN(n5282) );
  DFFRX1 \bArray_reg[12][31]  ( .D(n5898), .CK(clk), .RN(n7620), .Q(
        \bArray[12][31] ), .QN(n5093) );
  DFFRX1 \bArray_reg[12][30]  ( .D(n5897), .CK(clk), .RN(n7620), .Q(
        \bArray[12][30] ), .QN(n5092) );
  DFFRX1 \bArray_reg[12][29]  ( .D(n5896), .CK(clk), .RN(n7620), .Q(
        \bArray[12][29] ), .QN(n5091) );
  DFFRX1 \bArray_reg[12][28]  ( .D(n5895), .CK(clk), .RN(n7620), .Q(
        \bArray[12][28] ), .QN(n5090) );
  DFFRX1 \bArray_reg[2][31]  ( .D(n6378), .CK(clk), .RN(n7580), .Q(
        \bArray[2][31] ), .QN(n5573) );
  DFFRX1 \bArray_reg[2][30]  ( .D(n6377), .CK(clk), .RN(n7580), .Q(
        \bArray[2][30] ), .QN(n5572) );
  DFFRX1 \bArray_reg[2][29]  ( .D(n6376), .CK(clk), .RN(n7580), .Q(
        \bArray[2][29] ), .QN(n5571) );
  DFFRX1 \bArray_reg[2][28]  ( .D(n6375), .CK(clk), .RN(n7580), .Q(
        \bArray[2][28] ), .QN(n5570) );
  DFFRX1 \bArray_reg[6][31]  ( .D(n6186), .CK(clk), .RN(n7596), .Q(
        \bArray[6][31] ), .QN(n5381) );
  DFFRX1 \bArray_reg[6][30]  ( .D(n6185), .CK(clk), .RN(n7596), .Q(
        \bArray[6][30] ), .QN(n5380) );
  DFFRX1 \bArray_reg[6][29]  ( .D(n6184), .CK(clk), .RN(n7596), .Q(
        \bArray[6][29] ), .QN(n5379) );
  DFFRX1 \bArray_reg[6][28]  ( .D(n6183), .CK(clk), .RN(n7596), .Q(
        \bArray[6][28] ), .QN(n5378) );
  DFFRX1 \bArray_reg[10][31]  ( .D(n5994), .CK(clk), .RN(n7612), .Q(
        \bArray[10][31] ), .QN(n5189) );
  DFFRX1 \bArray_reg[10][30]  ( .D(n5993), .CK(clk), .RN(n7612), .Q(
        \bArray[10][30] ), .QN(n5188) );
  DFFRX1 \bArray_reg[10][29]  ( .D(n5992), .CK(clk), .RN(n7612), .Q(
        \bArray[10][29] ), .QN(n5187) );
  DFFRX1 \bArray_reg[10][28]  ( .D(n5991), .CK(clk), .RN(n7612), .Q(
        \bArray[10][28] ), .QN(n5186) );
  DFFRX1 \bArray_reg[14][31]  ( .D(n5802), .CK(clk), .RN(n7628), .Q(
        \bArray[14][31] ), .QN(n4997) );
  DFFRX1 \bArray_reg[14][30]  ( .D(n5801), .CK(clk), .RN(n7628), .Q(
        \bArray[14][30] ), .QN(n4996) );
  DFFRX1 \bArray_reg[14][29]  ( .D(n5800), .CK(clk), .RN(n7628), .Q(
        \bArray[14][29] ), .QN(n4995) );
  DFFRX1 \bArray_reg[14][28]  ( .D(n5799), .CK(clk), .RN(n7628), .Q(
        \bArray[14][28] ), .QN(n4994) );
  DFFQX1 \xArray_reg[1][34]  ( .D(N28739), .CK(clk), .Q(\xArray[1][34] ) );
  DFFQX1 \xArray_reg[1][33]  ( .D(N28738), .CK(clk), .Q(\xArray[1][33] ) );
  DFFQX1 \xArray_reg[13][34]  ( .D(N27971), .CK(clk), .Q(\xArray[13][34] ) );
  DFFQX1 \xArray_reg[13][33]  ( .D(N27970), .CK(clk), .Q(\xArray[13][33] ) );
  DFFQX1 \xArray_reg[9][34]  ( .D(N28227), .CK(clk), .Q(\xArray[9][34] ) );
  DFFQX1 \xArray_reg[9][33]  ( .D(N28226), .CK(clk), .Q(\xArray[9][33] ) );
  DFFQX1 \xArray_reg[8][34]  ( .D(N28291), .CK(clk), .Q(\xArray[8][34] ) );
  DFFQX1 \xArray_reg[8][33]  ( .D(N28290), .CK(clk), .Q(\xArray[8][33] ) );
  DFFQX1 \xArray_reg[10][34]  ( .D(N28163), .CK(clk), .Q(\xArray[10][34] ) );
  DFFQX1 \xArray_reg[10][33]  ( .D(N28162), .CK(clk), .Q(\xArray[10][33] ) );
  DFFQX1 \xArray_reg[6][34]  ( .D(N28419), .CK(clk), .Q(\xArray[6][34] ) );
  DFFQX1 \xArray_reg[6][33]  ( .D(N28418), .CK(clk), .Q(\xArray[6][33] ) );
  DFFQX1 \xArray_reg[15][31]  ( .D(N27840), .CK(clk), .Q(\xArray[15][31] ) );
  DFFQX1 \xArray_reg[5][31]  ( .D(N28480), .CK(clk), .Q(\xArray[5][31] ) );
  DFFQX1 \xArray_reg[4][31]  ( .D(N28544), .CK(clk), .Q(\xArray[4][31] ) );
  DFFQX1 \xArray_reg[14][31]  ( .D(N27904), .CK(clk), .Q(\xArray[14][31] ) );
  DFFQX1 \xArray_reg[11][31]  ( .D(N28096), .CK(clk), .Q(\xArray[11][31] ) );
  DFFQX1 \xArray_reg[1][32]  ( .D(N28737), .CK(clk), .Q(\xArray[1][32] ) );
  DFFQX1 \xArray_reg[7][31]  ( .D(N28352), .CK(clk), .Q(\xArray[7][31] ) );
  DFFQX1 \xArray_reg[13][32]  ( .D(N27969), .CK(clk), .Q(\xArray[13][32] ) );
  DFFQX1 \xArray_reg[9][32]  ( .D(N28225), .CK(clk), .Q(\xArray[9][32] ) );
  DFFQX1 \xArray_reg[8][32]  ( .D(N28289), .CK(clk), .Q(\xArray[8][32] ) );
  DFFQX1 \xArray_reg[10][32]  ( .D(N28161), .CK(clk), .Q(\xArray[10][32] ) );
  DFFQX1 \xArray_reg[6][32]  ( .D(N28417), .CK(clk), .Q(\xArray[6][32] ) );
  DFFQX1 \xArray_reg[9][31]  ( .D(N28224), .CK(clk), .Q(\xArray[9][31] ) );
  DFFQX1 \xArray_reg[8][31]  ( .D(N28288), .CK(clk), .Q(\xArray[8][31] ) );
  DFFRX1 \bArray_reg[1][27]  ( .D(n6422), .CK(clk), .RN(n7577), .Q(
        \bArray[1][27] ), .QN(n5617) );
  DFFRX1 \bArray_reg[1][26]  ( .D(n6421), .CK(clk), .RN(n7577), .Q(
        \bArray[1][26] ), .QN(n5616) );
  DFFRX1 \bArray_reg[5][27]  ( .D(n6230), .CK(clk), .RN(n7593), .Q(
        \bArray[5][27] ), .QN(n5425) );
  DFFRX1 \bArray_reg[5][26]  ( .D(n6229), .CK(clk), .RN(n7593), .Q(
        \bArray[5][26] ), .QN(n5424) );
  DFFRX1 \bArray_reg[9][27]  ( .D(n6038), .CK(clk), .RN(n7609), .Q(
        \bArray[9][27] ), .QN(n5233) );
  DFFRX1 \bArray_reg[9][26]  ( .D(n6037), .CK(clk), .RN(n7609), .Q(
        \bArray[9][26] ), .QN(n5232) );
  DFFRX1 \bArray_reg[13][27]  ( .D(n5846), .CK(clk), .RN(n7625), .Q(
        \bArray[13][27] ), .QN(n5041) );
  DFFRX1 \bArray_reg[13][26]  ( .D(n5845), .CK(clk), .RN(n7625), .Q(
        \bArray[13][26] ), .QN(n5040) );
  DFFRX1 \bArray_reg[3][27]  ( .D(n6326), .CK(clk), .RN(n7585), .Q(
        \bArray[3][27] ), .QN(n5521) );
  DFFRX1 \bArray_reg[3][26]  ( .D(n6325), .CK(clk), .RN(n7585), .Q(
        \bArray[3][26] ), .QN(n5520) );
  DFFRX1 \bArray_reg[7][27]  ( .D(n6134), .CK(clk), .RN(n7601), .Q(
        \bArray[7][27] ), .QN(n5329) );
  DFFRX1 \bArray_reg[7][26]  ( .D(n6133), .CK(clk), .RN(n7601), .Q(
        \bArray[7][26] ), .QN(n5328) );
  DFFRX1 \bArray_reg[11][27]  ( .D(n5942), .CK(clk), .RN(n7617), .Q(
        \bArray[11][27] ), .QN(n5137) );
  DFFRX1 \bArray_reg[11][26]  ( .D(n5941), .CK(clk), .RN(n7617), .Q(
        \bArray[11][26] ), .QN(n5136) );
  DFFRX1 \bArray_reg[15][27]  ( .D(n5750), .CK(clk), .RN(n7633), .Q(
        \bArray[15][27] ), .QN(n4945) );
  DFFRX1 \bArray_reg[15][26]  ( .D(n5749), .CK(clk), .RN(n7633), .Q(
        \bArray[15][26] ), .QN(n4944) );
  DFFRX1 \bArray_reg[0][27]  ( .D(n6470), .CK(clk), .RN(n7573), .Q(
        \bArray[0][27] ), .QN(n5665) );
  DFFRX1 \bArray_reg[0][26]  ( .D(n6469), .CK(clk), .RN(n7573), .Q(
        \bArray[0][26] ), .QN(n5664) );
  DFFRX1 \bArray_reg[4][27]  ( .D(n6278), .CK(clk), .RN(n7589), .Q(
        \bArray[4][27] ), .QN(n5473) );
  DFFRX1 \bArray_reg[4][26]  ( .D(n6277), .CK(clk), .RN(n7589), .Q(
        \bArray[4][26] ), .QN(n5472) );
  DFFRX1 \bArray_reg[8][27]  ( .D(n6086), .CK(clk), .RN(n7605), .Q(
        \bArray[8][27] ), .QN(n5281) );
  DFFRX1 \bArray_reg[8][26]  ( .D(n6085), .CK(clk), .RN(n7605), .Q(
        \bArray[8][26] ), .QN(n5280) );
  DFFRX1 \bArray_reg[12][27]  ( .D(n5894), .CK(clk), .RN(n7621), .Q(
        \bArray[12][27] ), .QN(n5089) );
  DFFRX1 \bArray_reg[12][26]  ( .D(n5893), .CK(clk), .RN(n7621), .Q(
        \bArray[12][26] ), .QN(n5088) );
  DFFRX1 \bArray_reg[2][27]  ( .D(n6374), .CK(clk), .RN(n7581), .Q(
        \bArray[2][27] ), .QN(n5569) );
  DFFRX1 \bArray_reg[2][26]  ( .D(n6373), .CK(clk), .RN(n7581), .Q(
        \bArray[2][26] ), .QN(n5568) );
  DFFRX1 \bArray_reg[6][27]  ( .D(n6182), .CK(clk), .RN(n7597), .Q(
        \bArray[6][27] ), .QN(n5377) );
  DFFRX1 \bArray_reg[6][26]  ( .D(n6181), .CK(clk), .RN(n7597), .Q(
        \bArray[6][26] ), .QN(n5376) );
  DFFRX1 \bArray_reg[10][27]  ( .D(n5990), .CK(clk), .RN(n7613), .Q(
        \bArray[10][27] ), .QN(n5185) );
  DFFRX1 \bArray_reg[10][26]  ( .D(n5989), .CK(clk), .RN(n7613), .Q(
        \bArray[10][26] ), .QN(n5184) );
  DFFRX1 \bArray_reg[14][27]  ( .D(n5798), .CK(clk), .RN(n7629), .Q(
        \bArray[14][27] ), .QN(n4993) );
  DFFRX1 \bArray_reg[14][26]  ( .D(n5797), .CK(clk), .RN(n7629), .Q(
        \bArray[14][26] ), .QN(n4992) );
  DFFQX1 \xArray_reg[15][30]  ( .D(N27839), .CK(clk), .Q(\xArray[15][30] ) );
  DFFQX1 \xArray_reg[15][29]  ( .D(N27838), .CK(clk), .Q(\xArray[15][29] ) );
  DFFQX1 \xArray_reg[0][31]  ( .D(N28800), .CK(clk), .Q(\xArray[0][31] ) );
  DFFQX1 \xArray_reg[0][30]  ( .D(N28799), .CK(clk), .Q(\xArray[0][30] ) );
  DFFQX1 \xArray_reg[5][30]  ( .D(N28479), .CK(clk), .Q(\xArray[5][30] ) );
  DFFQX1 \xArray_reg[5][29]  ( .D(N28478), .CK(clk), .Q(\xArray[5][29] ) );
  DFFQX1 \xArray_reg[4][30]  ( .D(N28543), .CK(clk), .Q(\xArray[4][30] ) );
  DFFQX1 \xArray_reg[14][30]  ( .D(N27903), .CK(clk), .Q(\xArray[14][30] ) );
  DFFQX1 \xArray_reg[11][30]  ( .D(N28095), .CK(clk), .Q(\xArray[11][30] ) );
  DFFQX1 \xArray_reg[11][29]  ( .D(N28094), .CK(clk), .Q(\xArray[11][29] ) );
  DFFQX1 \xArray_reg[12][31]  ( .D(N28032), .CK(clk), .Q(\xArray[12][31] ) );
  DFFQX1 \xArray_reg[12][30]  ( .D(N28031), .CK(clk), .Q(\xArray[12][30] ) );
  DFFQX1 \xArray_reg[7][30]  ( .D(N28351), .CK(clk), .Q(\xArray[7][30] ) );
  DFFQX1 \xArray_reg[7][29]  ( .D(N28350), .CK(clk), .Q(\xArray[7][29] ) );
  DFFQX1 \xArray_reg[1][31]  ( .D(N28736), .CK(clk), .Q(\xArray[1][31] ) );
  DFFQX1 \xArray_reg[1][30]  ( .D(N28735), .CK(clk), .Q(\xArray[1][30] ) );
  DFFQX1 \xArray_reg[13][31]  ( .D(N27968), .CK(clk), .Q(\xArray[13][31] ) );
  DFFQX1 \xArray_reg[13][30]  ( .D(N27967), .CK(clk), .Q(\xArray[13][30] ) );
  DFFQX1 \xArray_reg[9][30]  ( .D(N28223), .CK(clk), .Q(\xArray[9][30] ) );
  DFFQX1 \xArray_reg[8][30]  ( .D(N28287), .CK(clk), .Q(\xArray[8][30] ) );
  DFFQX1 \xArray_reg[15][28]  ( .D(N27837), .CK(clk), .Q(\xArray[15][28] ) );
  DFFQX1 \xArray_reg[15][27]  ( .D(N27836), .CK(clk), .Q(\xArray[15][27] ) );
  DFFQX1 \xArray_reg[0][29]  ( .D(N28798), .CK(clk), .Q(\xArray[0][29] ) );
  DFFQX1 \xArray_reg[0][28]  ( .D(N28797), .CK(clk), .Q(\xArray[0][28] ) );
  DFFQX1 \xArray_reg[5][28]  ( .D(N28477), .CK(clk), .Q(\xArray[5][28] ) );
  DFFQX1 \xArray_reg[5][27]  ( .D(N28476), .CK(clk), .Q(\xArray[5][27] ) );
  DFFQX1 \xArray_reg[4][29]  ( .D(N28542), .CK(clk), .Q(\xArray[4][29] ) );
  DFFQX1 \xArray_reg[4][28]  ( .D(N28541), .CK(clk), .Q(\xArray[4][28] ) );
  DFFQX1 \xArray_reg[11][28]  ( .D(N28093), .CK(clk), .Q(\xArray[11][28] ) );
  DFFQX1 \xArray_reg[11][27]  ( .D(N28092), .CK(clk), .Q(\xArray[11][27] ) );
  DFFQX1 \xArray_reg[12][29]  ( .D(N28030), .CK(clk), .Q(\xArray[12][29] ) );
  DFFQX1 \xArray_reg[12][28]  ( .D(N28029), .CK(clk), .Q(\xArray[12][28] ) );
  DFFQX1 \xArray_reg[7][28]  ( .D(N28349), .CK(clk), .Q(\xArray[7][28] ) );
  DFFQX1 \xArray_reg[7][27]  ( .D(N28348), .CK(clk), .Q(\xArray[7][27] ) );
  DFFQX1 \xArray_reg[1][29]  ( .D(N28734), .CK(clk), .Q(\xArray[1][29] ) );
  DFFQX1 \xArray_reg[1][28]  ( .D(N28733), .CK(clk), .Q(\xArray[1][28] ) );
  DFFQX1 \xArray_reg[13][29]  ( .D(N27966), .CK(clk), .Q(\xArray[13][29] ) );
  DFFQX1 \xArray_reg[13][28]  ( .D(N27965), .CK(clk), .Q(\xArray[13][28] ) );
  DFFQX1 \xArray_reg[9][29]  ( .D(N28222), .CK(clk), .Q(\xArray[9][29] ) );
  DFFQX1 \xArray_reg[8][29]  ( .D(N28286), .CK(clk), .Q(\xArray[8][29] ) );
  DFFQX1 \xArray_reg[8][28]  ( .D(N28285), .CK(clk), .Q(\xArray[8][28] ) );
  DFFQX1 \xArray_reg[15][26]  ( .D(N27835), .CK(clk), .Q(\xArray[15][26] ) );
  DFFQX1 \xArray_reg[15][25]  ( .D(N27834), .CK(clk), .Q(\xArray[15][25] ) );
  DFFQX1 \xArray_reg[0][27]  ( .D(N28796), .CK(clk), .Q(\xArray[0][27] ) );
  DFFQX1 \xArray_reg[0][26]  ( .D(N28795), .CK(clk), .Q(\xArray[0][26] ) );
  DFFQX1 \xArray_reg[5][26]  ( .D(N28475), .CK(clk), .Q(\xArray[5][26] ) );
  DFFQX1 \xArray_reg[5][25]  ( .D(N28474), .CK(clk), .Q(\xArray[5][25] ) );
  DFFQX1 \xArray_reg[4][27]  ( .D(N28540), .CK(clk), .Q(\xArray[4][27] ) );
  DFFQX1 \xArray_reg[4][26]  ( .D(N28539), .CK(clk), .Q(\xArray[4][26] ) );
  DFFQX1 \xArray_reg[11][26]  ( .D(N28091), .CK(clk), .Q(\xArray[11][26] ) );
  DFFQX1 \xArray_reg[11][25]  ( .D(N28090), .CK(clk), .Q(\xArray[11][25] ) );
  DFFQX1 \xArray_reg[12][27]  ( .D(N28028), .CK(clk), .Q(\xArray[12][27] ) );
  DFFQX1 \xArray_reg[12][26]  ( .D(N28027), .CK(clk), .Q(\xArray[12][26] ) );
  DFFQX1 \xArray_reg[7][26]  ( .D(N28347), .CK(clk), .Q(\xArray[7][26] ) );
  DFFQX1 \xArray_reg[7][25]  ( .D(N28346), .CK(clk), .Q(\xArray[7][25] ) );
  DFFQX1 \xArray_reg[1][27]  ( .D(N28732), .CK(clk), .Q(\xArray[1][27] ) );
  DFFQX1 \xArray_reg[1][26]  ( .D(N28731), .CK(clk), .Q(\xArray[1][26] ) );
  DFFQX1 \xArray_reg[13][27]  ( .D(N27964), .CK(clk), .Q(\xArray[13][27] ) );
  DFFQX1 \xArray_reg[13][26]  ( .D(N27963), .CK(clk), .Q(\xArray[13][26] ) );
  DFFQX1 \xArray_reg[8][27]  ( .D(N28284), .CK(clk), .Q(\xArray[8][27] ) );
  DFFQX1 \xArray_reg[8][26]  ( .D(N28283), .CK(clk), .Q(\xArray[8][26] ) );
  DFFQX1 \xArray_reg[3][24]  ( .D(N28601), .CK(clk), .Q(\xArray[3][24] ) );
  DFFQX1 \xArray_reg[0][25]  ( .D(N28794), .CK(clk), .Q(\xArray[0][25] ) );
  DFFQX1 \xArray_reg[5][24]  ( .D(N28473), .CK(clk), .Q(\xArray[5][24] ) );
  DFFQX1 \xArray_reg[4][25]  ( .D(N28538), .CK(clk), .Q(\xArray[4][25] ) );
  DFFQX1 \xArray_reg[12][25]  ( .D(N28026), .CK(clk), .Q(\xArray[12][25] ) );
  DFFQX1 \xArray_reg[7][24]  ( .D(N28345), .CK(clk), .Q(\xArray[7][24] ) );
  DFFQX1 \xArray_reg[1][25]  ( .D(N28730), .CK(clk), .Q(\xArray[1][25] ) );
  DFFQX1 \xArray_reg[13][25]  ( .D(N27962), .CK(clk), .Q(\xArray[13][25] ) );
  DFFRX1 \inCount_reg[1]  ( .D(N1807), .CK(clk), .RN(n7636), .Q(N1758), .QN(
        n5702) );
  DFFRX1 \inCount_reg[2]  ( .D(N1808), .CK(clk), .RN(n7636), .Q(N1759), .QN(
        n5703) );
  DFFRX1 \inCount_reg[3]  ( .D(N1809), .CK(clk), .RN(n7637), .Q(N1760), .QN(
        n74) );
  DFFRX1 \inCount_reg[0]  ( .D(N1806), .CK(clk), .RN(n7636), .Q(N1757), .QN(
        n5701) );
  DFFQX1 \xArray_reg[2][49]  ( .D(N28690), .CK(clk), .Q(\xArray[2][49] ) );
  DFFQX1 \xArray_reg[2][48]  ( .D(N28689), .CK(clk), .Q(\xArray[2][48] ) );
  DFFQX1 \xArray_reg[2][47]  ( .D(N28688), .CK(clk), .Q(\xArray[2][47] ) );
  DFFQX1 \xArray_reg[2][46]  ( .D(N28687), .CK(clk), .Q(\xArray[2][46] ) );
  DFFQX1 \xArray_reg[2][45]  ( .D(N28686), .CK(clk), .Q(\xArray[2][45] ) );
  DFFQX1 \xArray_reg[2][44]  ( .D(N28685), .CK(clk), .Q(\xArray[2][44] ) );
  DFFQX1 \xArray_reg[2][43]  ( .D(N28684), .CK(clk), .Q(\xArray[2][43] ) );
  DFFQX1 \xArray_reg[2][42]  ( .D(N28683), .CK(clk), .Q(\xArray[2][42] ) );
  DFFQX1 \xArray_reg[2][41]  ( .D(N28682), .CK(clk), .Q(\xArray[2][41] ) );
  DFFQX1 \xArray_reg[2][40]  ( .D(N28681), .CK(clk), .Q(\xArray[2][40] ) );
  DFFQX1 \xArray_reg[2][39]  ( .D(N28680), .CK(clk), .Q(\xArray[2][39] ) );
  DFFQX1 \xArray_reg[2][38]  ( .D(N28679), .CK(clk), .Q(\xArray[2][38] ) );
  DFFQX1 \xArray_reg[2][37]  ( .D(N28678), .CK(clk), .Q(\xArray[2][37] ) );
  DFFQX1 \xArray_reg[2][36]  ( .D(N28677), .CK(clk), .Q(\xArray[2][36] ) );
  DFFQX1 \xArray_reg[2][35]  ( .D(N28676), .CK(clk), .Q(\xArray[2][35] ) );
  DFFQX1 \xArray_reg[2][34]  ( .D(N28675), .CK(clk), .Q(\xArray[2][34] ) );
  DFFQX1 \xArray_reg[2][33]  ( .D(N28674), .CK(clk), .Q(\xArray[2][33] ) );
  DFFQX1 \xArray_reg[2][32]  ( .D(N28673), .CK(clk), .Q(\xArray[2][32] ) );
  DFFQX1 \xArray_reg[2][31]  ( .D(N28672), .CK(clk), .Q(\xArray[2][31] ) );
  DFFQX1 \xArray_reg[10][31]  ( .D(N28160), .CK(clk), .Q(\xArray[10][31] ) );
  DFFQX1 \xArray_reg[6][31]  ( .D(N28416), .CK(clk), .Q(\xArray[6][31] ) );
  DFFQX1 \xArray_reg[10][30]  ( .D(N28159), .CK(clk), .Q(\xArray[10][30] ) );
  DFFQX1 \xArray_reg[10][29]  ( .D(N28158), .CK(clk), .Q(\xArray[10][29] ) );
  DFFQX1 \xArray_reg[6][30]  ( .D(N28415), .CK(clk), .Q(\xArray[6][30] ) );
  DFFQX1 \xArray_reg[6][29]  ( .D(N28414), .CK(clk), .Q(\xArray[6][29] ) );
  DFFQX1 \xArray_reg[10][28]  ( .D(N28157), .CK(clk), .Q(\xArray[10][28] ) );
  DFFQX1 \xArray_reg[10][27]  ( .D(N28156), .CK(clk), .Q(\xArray[10][27] ) );
  DFFQX1 \xArray_reg[6][28]  ( .D(N28413), .CK(clk), .Q(\xArray[6][28] ) );
  DFFQX1 \xArray_reg[6][27]  ( .D(N28412), .CK(clk), .Q(\xArray[6][27] ) );
  DFFQX1 \xArray_reg[10][26]  ( .D(N28155), .CK(clk), .Q(\xArray[10][26] ) );
  DFFQX1 \xArray_reg[10][25]  ( .D(N28154), .CK(clk), .Q(\xArray[10][25] ) );
  DFFQX1 \xArray_reg[6][26]  ( .D(N28411), .CK(clk), .Q(\xArray[6][26] ) );
  DFFQX1 \xArray_reg[6][25]  ( .D(N28410), .CK(clk), .Q(\xArray[6][25] ) );
  DFFQX1 \xArray_reg[10][24]  ( .D(N28153), .CK(clk), .Q(\xArray[10][24] ) );
  DFFQXL \xArray_reg[15][41]  ( .D(N27850), .CK(clk), .Q(\xArray[15][41] ) );
  DFFQXL \xArray_reg[15][40]  ( .D(N27849), .CK(clk), .Q(\xArray[15][40] ) );
  DFFQXL \xArray_reg[14][41]  ( .D(N27914), .CK(clk), .Q(\xArray[14][41] ) );
  DFFQXL \xArray_reg[14][40]  ( .D(N27913), .CK(clk), .Q(\xArray[14][40] ) );
  DFFQXL \xArray_reg[0][41]  ( .D(N28810), .CK(clk), .Q(\xArray[0][41] ) );
  DFFQXL \xArray_reg[0][40]  ( .D(N28809), .CK(clk), .Q(\xArray[0][40] ) );
  DFFQXL \xArray_reg[11][41]  ( .D(N28106), .CK(clk), .Q(\xArray[11][41] ) );
  DFFQXL \xArray_reg[12][41]  ( .D(N28042), .CK(clk), .Q(\xArray[12][41] ) );
  DFFQXL \xArray_reg[11][40]  ( .D(N28105), .CK(clk), .Q(\xArray[11][40] ) );
  DFFQXL \xArray_reg[15][39]  ( .D(N27848), .CK(clk), .Q(\xArray[15][39] ) );
  DFFQXL \xArray_reg[14][39]  ( .D(N27912), .CK(clk), .Q(\xArray[14][39] ) );
  DFFQXL \xArray_reg[14][38]  ( .D(N27911), .CK(clk), .Q(\xArray[14][38] ) );
  DFFQXL \xArray_reg[0][39]  ( .D(N28808), .CK(clk), .Q(\xArray[0][39] ) );
  DFFQXL \xArray_reg[12][40]  ( .D(N28041), .CK(clk), .Q(\xArray[12][40] ) );
  DFFQXL \xArray_reg[15][37]  ( .D(N27846), .CK(clk), .Q(\xArray[15][37] ) );
  DFFQXL \xArray_reg[14][37]  ( .D(N27910), .CK(clk), .Q(\xArray[14][37] ) );
  DFFQXL \xArray_reg[14][36]  ( .D(N27909), .CK(clk), .Q(\xArray[14][36] ) );
  DFFQXL \xArray_reg[0][37]  ( .D(N28806), .CK(clk), .Q(\xArray[0][37] ) );
  DFFQXL \xArray_reg[15][36]  ( .D(N27845), .CK(clk), .Q(\xArray[15][36] ) );
  DFFQXL \xArray_reg[14][35]  ( .D(N27908), .CK(clk), .Q(\xArray[14][35] ) );
  DFFQXL \xArray_reg[0][36]  ( .D(N28805), .CK(clk), .Q(\xArray[0][36] ) );
  DFFQXL \xArray_reg[15][34]  ( .D(N27843), .CK(clk), .Q(\xArray[15][34] ) );
  DFFQXL \xArray_reg[15][33]  ( .D(N27842), .CK(clk), .Q(\xArray[15][33] ) );
  DFFQXL \xArray_reg[14][34]  ( .D(N27907), .CK(clk), .Q(\xArray[14][34] ) );
  DFFQXL \xArray_reg[14][33]  ( .D(N27906), .CK(clk), .Q(\xArray[14][33] ) );
  DFFQXL \xArray_reg[0][34]  ( .D(N28803), .CK(clk), .Q(\xArray[0][34] ) );
  DFFQXL \xArray_reg[0][33]  ( .D(N28802), .CK(clk), .Q(\xArray[0][33] ) );
  DFFQXL \xArray_reg[14][32]  ( .D(N27905), .CK(clk), .Q(\xArray[14][32] ) );
  DFFRX4 \xCount_reg[1]  ( .D(xCount_next[1]), .CK(clk), .RN(n7639), .Q(N1762), 
        .QN(n104) );
  DFFRX4 \xCount_reg[2]  ( .D(xCount_next[2]), .CK(clk), .RN(n7639), .Q(N1763), 
        .QN(n105) );
  DFFQX1 \xArray_reg[15][24]  ( .D(N27833), .CK(clk), .Q(\xArray[15][24] ) );
  DFFQX1 \xArray_reg[0][24]  ( .D(N28793), .CK(clk), .Q(\xArray[0][24] ) );
  DFFQX1 \xArray_reg[0][16]  ( .D(N28785), .CK(clk), .Q(\xArray[0][16] ) );
  DFFQX1 \xArray_reg[0][15]  ( .D(N28784), .CK(clk), .Q(\xArray[0][15] ) );
  DFFQX1 \xArray_reg[0][14]  ( .D(N28783), .CK(clk), .Q(\xArray[0][14] ) );
  DFFQX1 \xArray_reg[0][13]  ( .D(N28782), .CK(clk), .Q(\xArray[0][13] ) );
  DFFQX1 \xArray_reg[0][12]  ( .D(N28781), .CK(clk), .Q(\xArray[0][12] ) );
  DFFQX1 \xArray_reg[15][8]  ( .D(N27817), .CK(clk), .Q(\xArray[15][8] ) );
  DFFRX4 \xCount_reg[0]  ( .D(xCount_next[0]), .CK(clk), .RN(n7639), .Q(N1761), 
        .QN(n103) );
  DFFQXL \xArray_reg[3][63]  ( .D(N28640), .CK(clk), .Q(\xArray[3][63] ) );
  DFFQXL \xArray_reg[5][63]  ( .D(N28512), .CK(clk), .Q(\xArray[5][63] ) );
  DFFQXL \xArray_reg[4][63]  ( .D(N28576), .CK(clk), .Q(\xArray[4][63] ) );
  DFFQXL \xArray_reg[7][63]  ( .D(N28384), .CK(clk), .Q(\xArray[7][63] ) );
  DFFQXL \xArray_reg[15][63]  ( .D(N27872), .CK(clk), .Q(\xArray[15][63] ) );
  DFFQXL \xArray_reg[0][63]  ( .D(N28832), .CK(clk), .Q(\xArray[0][63] ) );
  DFFQXL \xArray_reg[11][63]  ( .D(N28128), .CK(clk), .Q(\xArray[11][63] ) );
  DFFQXL \xArray_reg[12][63]  ( .D(N28064), .CK(clk), .Q(\xArray[12][63] ) );
  DFFQXL \xArray_reg[3][62]  ( .D(N28639), .CK(clk), .Q(\xArray[3][62] ) );
  DFFQXL \xArray_reg[0][62]  ( .D(N28831), .CK(clk), .Q(\xArray[0][62] ) );
  DFFQXL \xArray_reg[4][62]  ( .D(N28575), .CK(clk), .Q(\xArray[4][62] ) );
  DFFQXL \xArray_reg[5][62]  ( .D(N28511), .CK(clk), .Q(\xArray[5][62] ) );
  DFFQXL \xArray_reg[12][62]  ( .D(N28063), .CK(clk), .Q(\xArray[12][62] ) );
  DFFQXL \xArray_reg[7][62]  ( .D(N28383), .CK(clk), .Q(\xArray[7][62] ) );
  DFFQXL \xArray_reg[3][61]  ( .D(N28638), .CK(clk), .Q(\xArray[3][61] ) );
  DFFQXL \xArray_reg[15][62]  ( .D(N27871), .CK(clk), .Q(\xArray[15][62] ) );
  DFFQXL \xArray_reg[4][61]  ( .D(N28574), .CK(clk), .Q(\xArray[4][61] ) );
  DFFQXL \xArray_reg[5][61]  ( .D(N28510), .CK(clk), .Q(\xArray[5][61] ) );
  DFFQXL \xArray_reg[11][62]  ( .D(N28127), .CK(clk), .Q(\xArray[11][62] ) );
  DFFQXL \xArray_reg[7][61]  ( .D(N28382), .CK(clk), .Q(\xArray[7][61] ) );
  DFFQXL \xArray_reg[3][60]  ( .D(N28637), .CK(clk), .Q(\xArray[3][60] ) );
  DFFQXL \xArray_reg[15][61]  ( .D(N27870), .CK(clk), .Q(\xArray[15][61] ) );
  DFFQXL \xArray_reg[0][61]  ( .D(N28830), .CK(clk), .Q(\xArray[0][61] ) );
  DFFQXL \xArray_reg[4][60]  ( .D(N28573), .CK(clk), .Q(\xArray[4][60] ) );
  DFFQXL \xArray_reg[5][60]  ( .D(N28509), .CK(clk), .Q(\xArray[5][60] ) );
  DFFQXL \xArray_reg[11][61]  ( .D(N28126), .CK(clk), .Q(\xArray[11][61] ) );
  DFFQXL \xArray_reg[12][61]  ( .D(N28062), .CK(clk), .Q(\xArray[12][61] ) );
  DFFQXL \xArray_reg[7][60]  ( .D(N28381), .CK(clk), .Q(\xArray[7][60] ) );
  DFFQXL \xArray_reg[3][59]  ( .D(N28636), .CK(clk), .Q(\xArray[3][59] ) );
  DFFQXL \xArray_reg[3][58]  ( .D(N28635), .CK(clk), .Q(\xArray[3][58] ) );
  DFFQXL \xArray_reg[15][60]  ( .D(N27869), .CK(clk), .Q(\xArray[15][60] ) );
  DFFQXL \xArray_reg[15][59]  ( .D(N27868), .CK(clk), .Q(\xArray[15][59] ) );
  DFFQXL \xArray_reg[15][58]  ( .D(N27867), .CK(clk), .Q(\xArray[15][58] ) );
  DFFQXL \xArray_reg[0][60]  ( .D(N28829), .CK(clk), .Q(\xArray[0][60] ) );
  DFFQXL \xArray_reg[0][59]  ( .D(N28828), .CK(clk), .Q(\xArray[0][59] ) );
  DFFQXL \xArray_reg[0][58]  ( .D(N28827), .CK(clk), .Q(\xArray[0][58] ) );
  DFFQXL \xArray_reg[4][59]  ( .D(N28572), .CK(clk), .Q(\xArray[4][59] ) );
  DFFQXL \xArray_reg[4][58]  ( .D(N28571), .CK(clk), .Q(\xArray[4][58] ) );
  DFFQXL \xArray_reg[5][59]  ( .D(N28508), .CK(clk), .Q(\xArray[5][59] ) );
  DFFQXL \xArray_reg[5][58]  ( .D(N28507), .CK(clk), .Q(\xArray[5][58] ) );
  DFFQXL \xArray_reg[11][60]  ( .D(N28125), .CK(clk), .Q(\xArray[11][60] ) );
  DFFQXL \xArray_reg[12][59]  ( .D(N28060), .CK(clk), .Q(\xArray[12][59] ) );
  DFFQXL \xArray_reg[12][58]  ( .D(N28059), .CK(clk), .Q(\xArray[12][58] ) );
  DFFQXL \xArray_reg[11][59]  ( .D(N28124), .CK(clk), .Q(\xArray[11][59] ) );
  DFFQXL \xArray_reg[11][58]  ( .D(N28123), .CK(clk), .Q(\xArray[11][58] ) );
  DFFQXL \xArray_reg[7][59]  ( .D(N28380), .CK(clk), .Q(\xArray[7][59] ) );
  DFFQXL \xArray_reg[7][58]  ( .D(N28379), .CK(clk), .Q(\xArray[7][58] ) );
  DFFQXL \xArray_reg[12][60]  ( .D(N28061), .CK(clk), .Q(\xArray[12][60] ) );
  DFFQXL \xArray_reg[3][57]  ( .D(N28634), .CK(clk), .Q(\xArray[3][57] ) );
  DFFQXL \xArray_reg[3][56]  ( .D(N28633), .CK(clk), .Q(\xArray[3][56] ) );
  DFFQXL \xArray_reg[15][57]  ( .D(N27866), .CK(clk), .Q(\xArray[15][57] ) );
  DFFQXL \xArray_reg[0][57]  ( .D(N28826), .CK(clk), .Q(\xArray[0][57] ) );
  DFFQXL \xArray_reg[4][56]  ( .D(N28569), .CK(clk), .Q(\xArray[4][56] ) );
  DFFQXL \xArray_reg[4][57]  ( .D(N28570), .CK(clk), .Q(\xArray[4][57] ) );
  DFFQXL \xArray_reg[5][57]  ( .D(N28506), .CK(clk), .Q(\xArray[5][57] ) );
  DFFQXL \xArray_reg[5][56]  ( .D(N28505), .CK(clk), .Q(\xArray[5][56] ) );
  DFFQXL \xArray_reg[12][57]  ( .D(N28058), .CK(clk), .Q(\xArray[12][57] ) );
  DFFQXL \xArray_reg[11][57]  ( .D(N28122), .CK(clk), .Q(\xArray[11][57] ) );
  DFFQXL \xArray_reg[7][56]  ( .D(N28377), .CK(clk), .Q(\xArray[7][56] ) );
  DFFQXL \xArray_reg[7][57]  ( .D(N28378), .CK(clk), .Q(\xArray[7][57] ) );
  DFFQXL \xArray_reg[3][55]  ( .D(N28632), .CK(clk), .Q(\xArray[3][55] ) );
  DFFQXL \xArray_reg[3][54]  ( .D(N28631), .CK(clk), .Q(\xArray[3][54] ) );
  DFFQXL \xArray_reg[15][55]  ( .D(N27864), .CK(clk), .Q(\xArray[15][55] ) );
  DFFQXL \xArray_reg[15][56]  ( .D(N27865), .CK(clk), .Q(\xArray[15][56] ) );
  DFFQXL \xArray_reg[0][56]  ( .D(N28825), .CK(clk), .Q(\xArray[0][56] ) );
  DFFQXL \xArray_reg[0][55]  ( .D(N28824), .CK(clk), .Q(\xArray[0][55] ) );
  DFFQXL \xArray_reg[5][54]  ( .D(N28503), .CK(clk), .Q(\xArray[5][54] ) );
  DFFQXL \xArray_reg[4][55]  ( .D(N28568), .CK(clk), .Q(\xArray[4][55] ) );
  DFFQXL \xArray_reg[4][54]  ( .D(N28567), .CK(clk), .Q(\xArray[4][54] ) );
  DFFQXL \xArray_reg[5][55]  ( .D(N28504), .CK(clk), .Q(\xArray[5][55] ) );
  DFFQXL \xArray_reg[12][56]  ( .D(N28057), .CK(clk), .Q(\xArray[12][56] ) );
  DFFQXL \xArray_reg[11][56]  ( .D(N28121), .CK(clk), .Q(\xArray[11][56] ) );
  DFFQXL \xArray_reg[12][55]  ( .D(N28056), .CK(clk), .Q(\xArray[12][55] ) );
  DFFQXL \xArray_reg[11][55]  ( .D(N28120), .CK(clk), .Q(\xArray[11][55] ) );
  DFFQXL \xArray_reg[7][55]  ( .D(N28376), .CK(clk), .Q(\xArray[7][55] ) );
  DFFQXL \xArray_reg[3][53]  ( .D(N28630), .CK(clk), .Q(\xArray[3][53] ) );
  DFFQXL \xArray_reg[15][54]  ( .D(N27863), .CK(clk), .Q(\xArray[15][54] ) );
  DFFQXL \xArray_reg[0][54]  ( .D(N28823), .CK(clk), .Q(\xArray[0][54] ) );
  DFFQXL \xArray_reg[5][53]  ( .D(N28502), .CK(clk), .Q(\xArray[5][53] ) );
  DFFQXL \xArray_reg[4][53]  ( .D(N28566), .CK(clk), .Q(\xArray[4][53] ) );
  DFFQXL \xArray_reg[12][54]  ( .D(N28055), .CK(clk), .Q(\xArray[12][54] ) );
  DFFQXL \xArray_reg[11][54]  ( .D(N28119), .CK(clk), .Q(\xArray[11][54] ) );
  DFFQXL \xArray_reg[7][54]  ( .D(N28375), .CK(clk), .Q(\xArray[7][54] ) );
  DFFQXL \xArray_reg[7][53]  ( .D(N28374), .CK(clk), .Q(\xArray[7][53] ) );
  DFFQXL \xArray_reg[3][52]  ( .D(N28629), .CK(clk), .Q(\xArray[3][52] ) );
  DFFQXL \xArray_reg[3][51]  ( .D(N28628), .CK(clk), .Q(\xArray[3][51] ) );
  DFFQXL \xArray_reg[15][53]  ( .D(N27862), .CK(clk), .Q(\xArray[15][53] ) );
  DFFQXL \xArray_reg[15][52]  ( .D(N27861), .CK(clk), .Q(\xArray[15][52] ) );
  DFFQXL \xArray_reg[0][53]  ( .D(N28822), .CK(clk), .Q(\xArray[0][53] ) );
  DFFQXL \xArray_reg[0][52]  ( .D(N28821), .CK(clk), .Q(\xArray[0][52] ) );
  DFFQXL \xArray_reg[5][52]  ( .D(N28501), .CK(clk), .Q(\xArray[5][52] ) );
  DFFQXL \xArray_reg[5][51]  ( .D(N28500), .CK(clk), .Q(\xArray[5][51] ) );
  DFFQXL \xArray_reg[4][52]  ( .D(N28565), .CK(clk), .Q(\xArray[4][52] ) );
  DFFQXL \xArray_reg[4][51]  ( .D(N28564), .CK(clk), .Q(\xArray[4][51] ) );
  DFFQXL \xArray_reg[12][53]  ( .D(N28054), .CK(clk), .Q(\xArray[12][53] ) );
  DFFQXL \xArray_reg[12][52]  ( .D(N28053), .CK(clk), .Q(\xArray[12][52] ) );
  DFFQXL \xArray_reg[11][53]  ( .D(N28118), .CK(clk), .Q(\xArray[11][53] ) );
  DFFQXL \xArray_reg[11][52]  ( .D(N28117), .CK(clk), .Q(\xArray[11][52] ) );
  DFFQXL \xArray_reg[7][52]  ( .D(N28373), .CK(clk), .Q(\xArray[7][52] ) );
  DFFQXL \xArray_reg[7][51]  ( .D(N28372), .CK(clk), .Q(\xArray[7][51] ) );
  DFFQXL \xArray_reg[3][50]  ( .D(N28627), .CK(clk), .Q(\xArray[3][50] ) );
  DFFQXL \xArray_reg[3][49]  ( .D(N28626), .CK(clk), .Q(\xArray[3][49] ) );
  DFFQXL \xArray_reg[15][50]  ( .D(N27859), .CK(clk), .Q(\xArray[15][50] ) );
  DFFQXL \xArray_reg[15][51]  ( .D(N27860), .CK(clk), .Q(\xArray[15][51] ) );
  DFFQXL \xArray_reg[0][51]  ( .D(N28820), .CK(clk), .Q(\xArray[0][51] ) );
  DFFQXL \xArray_reg[0][50]  ( .D(N28819), .CK(clk), .Q(\xArray[0][50] ) );
  DFFQXL \xArray_reg[5][50]  ( .D(N28499), .CK(clk), .Q(\xArray[5][50] ) );
  DFFQXL \xArray_reg[5][49]  ( .D(N28498), .CK(clk), .Q(\xArray[5][49] ) );
  DFFQXL \xArray_reg[4][50]  ( .D(N28563), .CK(clk), .Q(\xArray[4][50] ) );
  DFFQXL \xArray_reg[4][49]  ( .D(N28562), .CK(clk), .Q(\xArray[4][49] ) );
  DFFQXL \xArray_reg[12][51]  ( .D(N28052), .CK(clk), .Q(\xArray[12][51] ) );
  DFFQXL \xArray_reg[12][50]  ( .D(N28051), .CK(clk), .Q(\xArray[12][50] ) );
  DFFQXL \xArray_reg[11][50]  ( .D(N28115), .CK(clk), .Q(\xArray[11][50] ) );
  DFFQXL \xArray_reg[11][51]  ( .D(N28116), .CK(clk), .Q(\xArray[11][51] ) );
  DFFQXL \xArray_reg[7][50]  ( .D(N28371), .CK(clk), .Q(\xArray[7][50] ) );
  DFFQXL \xArray_reg[15][49]  ( .D(N27858), .CK(clk), .Q(\xArray[15][49] ) );
  DFFQXL \xArray_reg[14][49]  ( .D(N27922), .CK(clk), .Q(\xArray[14][49] ) );
  DFFQXL \xArray_reg[0][49]  ( .D(N28818), .CK(clk), .Q(\xArray[0][49] ) );
  DFFQXL \xArray_reg[12][49]  ( .D(N28050), .CK(clk), .Q(\xArray[12][49] ) );
  DFFQXL \xArray_reg[11][49]  ( .D(N28114), .CK(clk), .Q(\xArray[11][49] ) );
  DFFQXL \xArray_reg[7][49]  ( .D(N28370), .CK(clk), .Q(\xArray[7][49] ) );
  DFFQX1 \xArray_reg[7][41]  ( .D(N28362), .CK(clk), .Q(\xArray[7][41] ) );
  DFFQX1 \xArray_reg[7][40]  ( .D(N28361), .CK(clk), .Q(\xArray[7][40] ) );
  DFFQX1 \xArray_reg[7][39]  ( .D(N28360), .CK(clk), .Q(\xArray[7][39] ) );
  DFFQX1 \xArray_reg[0][38]  ( .D(N28807), .CK(clk), .Q(\xArray[0][38] ) );
  DFFQX1 \xArray_reg[11][39]  ( .D(N28104), .CK(clk), .Q(\xArray[11][39] ) );
  DFFQX1 \xArray_reg[12][39]  ( .D(N28040), .CK(clk), .Q(\xArray[12][39] ) );
  DFFQX1 \xArray_reg[11][38]  ( .D(N28103), .CK(clk), .Q(\xArray[11][38] ) );
  DFFQX1 \xArray_reg[12][38]  ( .D(N28039), .CK(clk), .Q(\xArray[12][38] ) );
  DFFQX1 \xArray_reg[7][38]  ( .D(N28359), .CK(clk), .Q(\xArray[7][38] ) );
  DFFQX1 \xArray_reg[7][37]  ( .D(N28358), .CK(clk), .Q(\xArray[7][37] ) );
  DFFQX1 \xArray_reg[11][37]  ( .D(N28102), .CK(clk), .Q(\xArray[11][37] ) );
  DFFQX1 \xArray_reg[12][37]  ( .D(N28038), .CK(clk), .Q(\xArray[12][37] ) );
  DFFQX1 \xArray_reg[11][36]  ( .D(N28101), .CK(clk), .Q(\xArray[11][36] ) );
  DFFQX1 \xArray_reg[12][36]  ( .D(N28037), .CK(clk), .Q(\xArray[12][36] ) );
  DFFQX1 \xArray_reg[7][36]  ( .D(N28357), .CK(clk), .Q(\xArray[7][36] ) );
  DFFQX1 \xArray_reg[7][35]  ( .D(N28356), .CK(clk), .Q(\xArray[7][35] ) );
  DFFQX1 \xArray_reg[0][35]  ( .D(N28804), .CK(clk), .Q(\xArray[0][35] ) );
  DFFQX1 \xArray_reg[11][34]  ( .D(N28099), .CK(clk), .Q(\xArray[11][34] ) );
  DFFQX1 \xArray_reg[12][34]  ( .D(N28035), .CK(clk), .Q(\xArray[12][34] ) );
  DFFQX1 \xArray_reg[11][35]  ( .D(N28100), .CK(clk), .Q(\xArray[11][35] ) );
  DFFQX1 \xArray_reg[12][35]  ( .D(N28036), .CK(clk), .Q(\xArray[12][35] ) );
  DFFQX1 \xArray_reg[7][34]  ( .D(N28355), .CK(clk), .Q(\xArray[7][34] ) );
  DFFQX1 \xArray_reg[7][33]  ( .D(N28354), .CK(clk), .Q(\xArray[7][33] ) );
  DFFQX1 \xArray_reg[11][33]  ( .D(N28098), .CK(clk), .Q(\xArray[11][33] ) );
  DFFQX1 \xArray_reg[12][33]  ( .D(N28034), .CK(clk), .Q(\xArray[12][33] ) );
  DFFQX1 \xArray_reg[9][28]  ( .D(N28221), .CK(clk), .Q(\xArray[9][28] ) );
  DFFQX1 \xArray_reg[4][24]  ( .D(N28537), .CK(clk), .Q(\xArray[4][24] ) );
  DFFQX1 \xArray_reg[11][24]  ( .D(N28089), .CK(clk), .Q(\xArray[11][24] ) );
  DFFQX1 \xArray_reg[12][24]  ( .D(N28025), .CK(clk), .Q(\xArray[12][24] ) );
  DFFQX1 \xArray_reg[8][25]  ( .D(N28282), .CK(clk), .Q(\xArray[8][25] ) );
  DFFQXL \xArray_reg[4][41]  ( .D(N28554), .CK(clk), .Q(\xArray[4][41] ) );
  DFFQXL \xArray_reg[5][41]  ( .D(N28490), .CK(clk), .Q(\xArray[5][41] ) );
  DFFQXL \xArray_reg[5][40]  ( .D(N28489), .CK(clk), .Q(\xArray[5][40] ) );
  DFFQXL \xArray_reg[3][41]  ( .D(N28618), .CK(clk), .Q(\xArray[3][41] ) );
  DFFQXL \xArray_reg[3][40]  ( .D(N28617), .CK(clk), .Q(\xArray[3][40] ) );
  DFFQXL \xArray_reg[4][40]  ( .D(N28553), .CK(clk), .Q(\xArray[4][40] ) );
  DFFQXL \xArray_reg[4][39]  ( .D(N28552), .CK(clk), .Q(\xArray[4][39] ) );
  DFFQXL \xArray_reg[5][39]  ( .D(N28488), .CK(clk), .Q(\xArray[5][39] ) );
  DFFQXL \xArray_reg[3][38]  ( .D(N28615), .CK(clk), .Q(\xArray[3][38] ) );
  DFFQXL \xArray_reg[3][39]  ( .D(N28616), .CK(clk), .Q(\xArray[3][39] ) );
  DFFQXL \xArray_reg[15][38]  ( .D(N27847), .CK(clk), .Q(\xArray[15][38] ) );
  DFFQXL \xArray_reg[4][37]  ( .D(N28550), .CK(clk), .Q(\xArray[4][37] ) );
  DFFQXL \xArray_reg[4][38]  ( .D(N28551), .CK(clk), .Q(\xArray[4][38] ) );
  DFFQXL \xArray_reg[5][38]  ( .D(N28487), .CK(clk), .Q(\xArray[5][38] ) );
  DFFQXL \xArray_reg[5][37]  ( .D(N28486), .CK(clk), .Q(\xArray[5][37] ) );
  DFFQXL \xArray_reg[3][36]  ( .D(N28613), .CK(clk), .Q(\xArray[3][36] ) );
  DFFQXL \xArray_reg[3][37]  ( .D(N28614), .CK(clk), .Q(\xArray[3][37] ) );
  DFFQXL \xArray_reg[15][35]  ( .D(N27844), .CK(clk), .Q(\xArray[15][35] ) );
  DFFQXL \xArray_reg[4][36]  ( .D(N28549), .CK(clk), .Q(\xArray[4][36] ) );
  DFFQXL \xArray_reg[4][35]  ( .D(N28548), .CK(clk), .Q(\xArray[4][35] ) );
  DFFQXL \xArray_reg[5][36]  ( .D(N28485), .CK(clk), .Q(\xArray[5][36] ) );
  DFFQXL \xArray_reg[5][35]  ( .D(N28484), .CK(clk), .Q(\xArray[5][35] ) );
  DFFQXL \xArray_reg[3][35]  ( .D(N28612), .CK(clk), .Q(\xArray[3][35] ) );
  DFFQXL \xArray_reg[4][34]  ( .D(N28547), .CK(clk), .Q(\xArray[4][34] ) );
  DFFQXL \xArray_reg[5][33]  ( .D(N28482), .CK(clk), .Q(\xArray[5][33] ) );
  DFFQXL \xArray_reg[5][34]  ( .D(N28483), .CK(clk), .Q(\xArray[5][34] ) );
  DFFQX1 \xArray_reg[2][55]  ( .D(N28696), .CK(clk), .Q(\xArray[2][55] ) );
  DFFQX1 \xArray_reg[2][54]  ( .D(N28695), .CK(clk), .Q(\xArray[2][54] ) );
  DFFQX1 \xArray_reg[2][53]  ( .D(N28694), .CK(clk), .Q(\xArray[2][53] ) );
  DFFQX1 \xArray_reg[2][52]  ( .D(N28693), .CK(clk), .Q(\xArray[2][52] ) );
  DFFQX1 \xArray_reg[2][51]  ( .D(N28692), .CK(clk), .Q(\xArray[2][51] ) );
  DFFQX1 \xArray_reg[2][50]  ( .D(N28691), .CK(clk), .Q(\xArray[2][50] ) );
  DFFRX1 \bArray_reg[2][24]  ( .D(n6371), .CK(clk), .RN(n7581), .Q(
        \bArray[2][24] ), .QN(n5566) );
  DFFRX1 \bArray_reg[6][24]  ( .D(n6179), .CK(clk), .RN(n7597), .Q(
        \bArray[6][24] ), .QN(n5374) );
  DFFRX1 \bArray_reg[10][24]  ( .D(n5987), .CK(clk), .RN(n7613), .Q(
        \bArray[10][24] ), .QN(n5182) );
  DFFRX1 \bArray_reg[14][24]  ( .D(n5795), .CK(clk), .RN(n7629), .Q(
        \bArray[14][24] ), .QN(n4990) );
  DFFRX1 \bArray_reg[1][24]  ( .D(n6419), .CK(clk), .RN(n7577), .Q(
        \bArray[1][24] ), .QN(n5614) );
  DFFRX1 \bArray_reg[5][24]  ( .D(n6227), .CK(clk), .RN(n7593), .Q(
        \bArray[5][24] ), .QN(n5422) );
  DFFRX1 \bArray_reg[9][24]  ( .D(n6035), .CK(clk), .RN(n7609), .Q(
        \bArray[9][24] ), .QN(n5230) );
  DFFRX1 \bArray_reg[13][24]  ( .D(n5843), .CK(clk), .RN(n7625), .Q(
        \bArray[13][24] ), .QN(n5038) );
  DFFRX1 \bArray_reg[3][24]  ( .D(n6323), .CK(clk), .RN(n7585), .Q(
        \bArray[3][24] ), .QN(n5518) );
  DFFRX1 \bArray_reg[7][24]  ( .D(n6131), .CK(clk), .RN(n7601), .Q(
        \bArray[7][24] ), .QN(n5326) );
  DFFRX1 \bArray_reg[11][24]  ( .D(n5939), .CK(clk), .RN(n7617), .Q(
        \bArray[11][24] ), .QN(n5134) );
  DFFRX1 \bArray_reg[15][24]  ( .D(n5747), .CK(clk), .RN(n7633), .Q(
        \bArray[15][24] ), .QN(n4942) );
  DFFRX1 \bArray_reg[0][24]  ( .D(n6467), .CK(clk), .RN(n7573), .Q(
        \bArray[0][24] ), .QN(n5662) );
  DFFRX1 \bArray_reg[4][24]  ( .D(n6275), .CK(clk), .RN(n7589), .Q(
        \bArray[4][24] ), .QN(n5470) );
  DFFRX1 \bArray_reg[8][24]  ( .D(n6083), .CK(clk), .RN(n7605), .Q(
        \bArray[8][24] ), .QN(n5278) );
  DFFRX1 \bArray_reg[12][24]  ( .D(n5891), .CK(clk), .RN(n7621), .Q(
        \bArray[12][24] ), .QN(n5086) );
  DFFRX1 \bArray_reg[2][25]  ( .D(n6372), .CK(clk), .RN(n7581), .Q(
        \bArray[2][25] ), .QN(n5567) );
  DFFRX1 \bArray_reg[6][25]  ( .D(n6180), .CK(clk), .RN(n7597), .Q(
        \bArray[6][25] ), .QN(n5375) );
  DFFRX1 \bArray_reg[10][25]  ( .D(n5988), .CK(clk), .RN(n7613), .Q(
        \bArray[10][25] ), .QN(n5183) );
  DFFRX1 \bArray_reg[14][25]  ( .D(n5796), .CK(clk), .RN(n7629), .Q(
        \bArray[14][25] ), .QN(n4991) );
  DFFRX1 \bArray_reg[1][25]  ( .D(n6420), .CK(clk), .RN(n7577), .Q(
        \bArray[1][25] ), .QN(n5615) );
  DFFRX1 \bArray_reg[5][25]  ( .D(n6228), .CK(clk), .RN(n7593), .Q(
        \bArray[5][25] ), .QN(n5423) );
  DFFRX1 \bArray_reg[9][25]  ( .D(n6036), .CK(clk), .RN(n7609), .Q(
        \bArray[9][25] ), .QN(n5231) );
  DFFRX1 \bArray_reg[13][25]  ( .D(n5844), .CK(clk), .RN(n7625), .Q(
        \bArray[13][25] ), .QN(n5039) );
  DFFRX1 \bArray_reg[3][25]  ( .D(n6324), .CK(clk), .RN(n7585), .Q(
        \bArray[3][25] ), .QN(n5519) );
  DFFRX1 \bArray_reg[7][25]  ( .D(n6132), .CK(clk), .RN(n7601), .Q(
        \bArray[7][25] ), .QN(n5327) );
  DFFRX1 \bArray_reg[11][25]  ( .D(n5940), .CK(clk), .RN(n7617), .Q(
        \bArray[11][25] ), .QN(n5135) );
  DFFRX1 \bArray_reg[15][25]  ( .D(n5748), .CK(clk), .RN(n7633), .Q(
        \bArray[15][25] ), .QN(n4943) );
  DFFRX1 \bArray_reg[0][25]  ( .D(n6468), .CK(clk), .RN(n7573), .Q(
        \bArray[0][25] ), .QN(n5663) );
  DFFRX1 \bArray_reg[4][25]  ( .D(n6276), .CK(clk), .RN(n7589), .Q(
        \bArray[4][25] ), .QN(n5471) );
  DFFRX1 \bArray_reg[8][25]  ( .D(n6084), .CK(clk), .RN(n7605), .Q(
        \bArray[8][25] ), .QN(n5279) );
  DFFRX1 \bArray_reg[12][25]  ( .D(n5892), .CK(clk), .RN(n7621), .Q(
        \bArray[12][25] ), .QN(n5087) );
  DFFRX1 \bArray_reg[2][23]  ( .D(n6370), .CK(clk), .RN(n7581), .Q(
        \bArray[2][23] ), .QN(n5565) );
  DFFRX1 \bArray_reg[6][23]  ( .D(n6178), .CK(clk), .RN(n7597), .Q(
        \bArray[6][23] ), .QN(n5373) );
  DFFRX1 \bArray_reg[10][23]  ( .D(n5986), .CK(clk), .RN(n7613), .Q(
        \bArray[10][23] ), .QN(n5181) );
  DFFRX1 \bArray_reg[14][23]  ( .D(n5794), .CK(clk), .RN(n7629), .Q(
        \bArray[14][23] ), .QN(n4989) );
  DFFRX1 \bArray_reg[1][23]  ( .D(n6418), .CK(clk), .RN(n7577), .Q(
        \bArray[1][23] ), .QN(n5613) );
  DFFRX1 \bArray_reg[1][22]  ( .D(n6417), .CK(clk), .RN(n7577), .Q(
        \bArray[1][22] ), .QN(n5612) );
  DFFRX1 \bArray_reg[5][23]  ( .D(n6226), .CK(clk), .RN(n7593), .Q(
        \bArray[5][23] ), .QN(n5421) );
  DFFRX1 \bArray_reg[9][23]  ( .D(n6034), .CK(clk), .RN(n7609), .Q(
        \bArray[9][23] ), .QN(n5229) );
  DFFRX1 \bArray_reg[13][23]  ( .D(n5842), .CK(clk), .RN(n7625), .Q(
        \bArray[13][23] ), .QN(n5037) );
  DFFRX1 \bArray_reg[3][23]  ( .D(n6322), .CK(clk), .RN(n7585), .Q(
        \bArray[3][23] ), .QN(n5517) );
  DFFRX1 \bArray_reg[7][23]  ( .D(n6130), .CK(clk), .RN(n7601), .Q(
        \bArray[7][23] ), .QN(n5325) );
  DFFRX1 \bArray_reg[11][23]  ( .D(n5938), .CK(clk), .RN(n7617), .Q(
        \bArray[11][23] ), .QN(n5133) );
  DFFRX1 \bArray_reg[15][23]  ( .D(n5746), .CK(clk), .RN(n7633), .Q(
        \bArray[15][23] ), .QN(n4941) );
  DFFRX1 \bArray_reg[0][23]  ( .D(n6466), .CK(clk), .RN(n7573), .Q(
        \bArray[0][23] ), .QN(n5661) );
  DFFRX1 \bArray_reg[0][22]  ( .D(n6465), .CK(clk), .RN(n7573), .Q(
        \bArray[0][22] ), .QN(n5660) );
  DFFRX1 \bArray_reg[4][23]  ( .D(n6274), .CK(clk), .RN(n7589), .Q(
        \bArray[4][23] ), .QN(n5469) );
  DFFRX1 \bArray_reg[8][23]  ( .D(n6082), .CK(clk), .RN(n7605), .Q(
        \bArray[8][23] ), .QN(n5277) );
  DFFRX1 \bArray_reg[12][23]  ( .D(n5890), .CK(clk), .RN(n7621), .Q(
        \bArray[12][23] ), .QN(n5085) );
  DFFRX1 \bArray_reg[6][22]  ( .D(n6177), .CK(clk), .RN(n7597), .Q(
        \bArray[6][22] ), .QN(n5372) );
  DFFRX1 \bArray_reg[10][22]  ( .D(n5985), .CK(clk), .RN(n7613), .Q(
        \bArray[10][22] ), .QN(n5180) );
  DFFRX1 \bArray_reg[14][22]  ( .D(n5793), .CK(clk), .RN(n7629), .Q(
        \bArray[14][22] ), .QN(n4988) );
  DFFRX1 \bArray_reg[5][22]  ( .D(n6225), .CK(clk), .RN(n7593), .Q(
        \bArray[5][22] ), .QN(n5420) );
  DFFRX1 \bArray_reg[9][22]  ( .D(n6033), .CK(clk), .RN(n7609), .Q(
        \bArray[9][22] ), .QN(n5228) );
  DFFRX1 \bArray_reg[13][22]  ( .D(n5841), .CK(clk), .RN(n7625), .Q(
        \bArray[13][22] ), .QN(n5036) );
  DFFRX1 \bArray_reg[7][22]  ( .D(n6129), .CK(clk), .RN(n7601), .Q(
        \bArray[7][22] ), .QN(n5324) );
  DFFRX1 \bArray_reg[11][22]  ( .D(n5937), .CK(clk), .RN(n7617), .Q(
        \bArray[11][22] ), .QN(n5132) );
  DFFRX1 \bArray_reg[15][22]  ( .D(n5745), .CK(clk), .RN(n7633), .Q(
        \bArray[15][22] ), .QN(n4940) );
  DFFRX1 \bArray_reg[4][22]  ( .D(n6273), .CK(clk), .RN(n7589), .Q(
        \bArray[4][22] ), .QN(n5468) );
  DFFRX1 \bArray_reg[8][22]  ( .D(n6081), .CK(clk), .RN(n7605), .Q(
        \bArray[8][22] ), .QN(n5276) );
  DFFRX1 \bArray_reg[12][22]  ( .D(n5889), .CK(clk), .RN(n7621), .Q(
        \bArray[12][22] ), .QN(n5084) );
  DFFRX1 \bArray_reg[2][22]  ( .D(n6369), .CK(clk), .RN(n7581), .Q(
        \bArray[2][22] ), .QN(n5564) );
  DFFRX1 \bArray_reg[6][21]  ( .D(n6176), .CK(clk), .RN(n7597), .Q(
        \bArray[6][21] ), .QN(n5371) );
  DFFRX1 \bArray_reg[10][21]  ( .D(n5984), .CK(clk), .RN(n7613), .Q(
        \bArray[10][21] ), .QN(n5179) );
  DFFRX1 \bArray_reg[14][21]  ( .D(n5792), .CK(clk), .RN(n7629), .Q(
        \bArray[14][21] ), .QN(n4987) );
  DFFRX1 \bArray_reg[5][21]  ( .D(n6224), .CK(clk), .RN(n7593), .Q(
        \bArray[5][21] ), .QN(n5419) );
  DFFRX1 \bArray_reg[9][21]  ( .D(n6032), .CK(clk), .RN(n7609), .Q(
        \bArray[9][21] ), .QN(n5227) );
  DFFRX1 \bArray_reg[13][21]  ( .D(n5840), .CK(clk), .RN(n7625), .Q(
        \bArray[13][21] ), .QN(n5035) );
  DFFRX1 \bArray_reg[3][22]  ( .D(n6321), .CK(clk), .RN(n7585), .Q(
        \bArray[3][22] ), .QN(n5516) );
  DFFRX1 \bArray_reg[7][21]  ( .D(n6128), .CK(clk), .RN(n7601), .Q(
        \bArray[7][21] ), .QN(n5323) );
  DFFRX1 \bArray_reg[11][21]  ( .D(n5936), .CK(clk), .RN(n7617), .Q(
        \bArray[11][21] ), .QN(n5131) );
  DFFRX1 \bArray_reg[15][21]  ( .D(n5744), .CK(clk), .RN(n7633), .Q(
        \bArray[15][21] ), .QN(n4939) );
  DFFRX1 \bArray_reg[4][21]  ( .D(n6272), .CK(clk), .RN(n7589), .Q(
        \bArray[4][21] ), .QN(n5467) );
  DFFRX1 \bArray_reg[8][21]  ( .D(n6080), .CK(clk), .RN(n7605), .Q(
        \bArray[8][21] ), .QN(n5275) );
  DFFRX1 \bArray_reg[12][21]  ( .D(n5888), .CK(clk), .RN(n7621), .Q(
        \bArray[12][21] ), .QN(n5083) );
  DFFRX1 \bArray_reg[2][21]  ( .D(n6368), .CK(clk), .RN(n7581), .Q(
        \bArray[2][21] ), .QN(n5563) );
  DFFRX1 \bArray_reg[1][21]  ( .D(n6416), .CK(clk), .RN(n7577), .Q(
        \bArray[1][21] ), .QN(n5611) );
  DFFRX1 \bArray_reg[3][21]  ( .D(n6320), .CK(clk), .RN(n7585), .Q(
        \bArray[3][21] ), .QN(n5515) );
  DFFRX1 \bArray_reg[0][21]  ( .D(n6464), .CK(clk), .RN(n7573), .Q(
        \bArray[0][21] ), .QN(n5659) );
  DFFRX1 \bArray_reg[2][20]  ( .D(n6367), .CK(clk), .RN(n7581), .Q(
        \bArray[2][20] ), .QN(n5562) );
  DFFRX1 \bArray_reg[2][19]  ( .D(n6366), .CK(clk), .RN(n7581), .Q(
        \bArray[2][19] ), .QN(n5561) );
  DFFRX1 \bArray_reg[6][20]  ( .D(n6175), .CK(clk), .RN(n7597), .Q(
        \bArray[6][20] ), .QN(n5370) );
  DFFRX1 \bArray_reg[6][19]  ( .D(n6174), .CK(clk), .RN(n7597), .Q(
        \bArray[6][19] ), .QN(n5369) );
  DFFRX1 \bArray_reg[10][20]  ( .D(n5983), .CK(clk), .RN(n7613), .Q(
        \bArray[10][20] ), .QN(n5178) );
  DFFRX1 \bArray_reg[10][19]  ( .D(n5982), .CK(clk), .RN(n7613), .Q(
        \bArray[10][19] ), .QN(n5177) );
  DFFRX1 \bArray_reg[14][20]  ( .D(n5791), .CK(clk), .RN(n7629), .Q(
        \bArray[14][20] ), .QN(n4986) );
  DFFRX1 \bArray_reg[14][19]  ( .D(n5790), .CK(clk), .RN(n7629), .Q(
        \bArray[14][19] ), .QN(n4985) );
  DFFRX1 \bArray_reg[1][20]  ( .D(n6415), .CK(clk), .RN(n7577), .Q(
        \bArray[1][20] ), .QN(n5610) );
  DFFRX1 \bArray_reg[1][19]  ( .D(n6414), .CK(clk), .RN(n7577), .Q(
        \bArray[1][19] ), .QN(n5609) );
  DFFRX1 \bArray_reg[5][20]  ( .D(n6223), .CK(clk), .RN(n7593), .Q(
        \bArray[5][20] ), .QN(n5418) );
  DFFRX1 \bArray_reg[5][19]  ( .D(n6222), .CK(clk), .RN(n7593), .Q(
        \bArray[5][19] ), .QN(n5417) );
  DFFRX1 \bArray_reg[9][20]  ( .D(n6031), .CK(clk), .RN(n7609), .Q(
        \bArray[9][20] ), .QN(n5226) );
  DFFRX1 \bArray_reg[9][19]  ( .D(n6030), .CK(clk), .RN(n7609), .Q(
        \bArray[9][19] ), .QN(n5225) );
  DFFRX1 \bArray_reg[13][20]  ( .D(n5839), .CK(clk), .RN(n7625), .Q(
        \bArray[13][20] ), .QN(n5034) );
  DFFRX1 \bArray_reg[13][19]  ( .D(n5838), .CK(clk), .RN(n7625), .Q(
        \bArray[13][19] ), .QN(n5033) );
  DFFRX1 \bArray_reg[3][20]  ( .D(n6319), .CK(clk), .RN(n7585), .Q(
        \bArray[3][20] ), .QN(n5514) );
  DFFRX1 \bArray_reg[3][19]  ( .D(n6318), .CK(clk), .RN(n7585), .Q(
        \bArray[3][19] ), .QN(n5513) );
  DFFRX1 \bArray_reg[7][20]  ( .D(n6127), .CK(clk), .RN(n7601), .Q(
        \bArray[7][20] ), .QN(n5322) );
  DFFRX1 \bArray_reg[7][19]  ( .D(n6126), .CK(clk), .RN(n7601), .Q(
        \bArray[7][19] ), .QN(n5321) );
  DFFRX1 \bArray_reg[11][20]  ( .D(n5935), .CK(clk), .RN(n7617), .Q(
        \bArray[11][20] ), .QN(n5130) );
  DFFRX1 \bArray_reg[11][19]  ( .D(n5934), .CK(clk), .RN(n7617), .Q(
        \bArray[11][19] ), .QN(n5129) );
  DFFRX1 \bArray_reg[15][20]  ( .D(n5743), .CK(clk), .RN(n7633), .Q(
        \bArray[15][20] ), .QN(n4938) );
  DFFRX1 \bArray_reg[15][19]  ( .D(n5742), .CK(clk), .RN(n7633), .Q(
        \bArray[15][19] ), .QN(n4937) );
  DFFRX1 \bArray_reg[0][20]  ( .D(n6463), .CK(clk), .RN(n7573), .Q(
        \bArray[0][20] ), .QN(n5658) );
  DFFRX1 \bArray_reg[0][19]  ( .D(n6462), .CK(clk), .RN(n7573), .Q(
        \bArray[0][19] ), .QN(n5657) );
  DFFRX1 \bArray_reg[4][20]  ( .D(n6271), .CK(clk), .RN(n7589), .Q(
        \bArray[4][20] ), .QN(n5466) );
  DFFRX1 \bArray_reg[4][19]  ( .D(n6270), .CK(clk), .RN(n7589), .Q(
        \bArray[4][19] ), .QN(n5465) );
  DFFRX1 \bArray_reg[8][20]  ( .D(n6079), .CK(clk), .RN(n7605), .Q(
        \bArray[8][20] ), .QN(n5274) );
  DFFRX1 \bArray_reg[8][19]  ( .D(n6078), .CK(clk), .RN(n7605), .Q(
        \bArray[8][19] ), .QN(n5273) );
  DFFRX1 \bArray_reg[12][20]  ( .D(n5887), .CK(clk), .RN(n7621), .Q(
        \bArray[12][20] ), .QN(n5082) );
  DFFRX1 \bArray_reg[12][19]  ( .D(n5886), .CK(clk), .RN(n7621), .Q(
        \bArray[12][19] ), .QN(n5081) );
  DFFRX1 \bArray_reg[2][18]  ( .D(n6365), .CK(clk), .RN(n7581), .Q(
        \bArray[2][18] ), .QN(n5560) );
  DFFRX1 \bArray_reg[6][18]  ( .D(n6173), .CK(clk), .RN(n7597), .Q(
        \bArray[6][18] ), .QN(n5368) );
  DFFRX1 \bArray_reg[1][18]  ( .D(n6413), .CK(clk), .RN(n7577), .Q(
        \bArray[1][18] ), .QN(n5608) );
  DFFRX1 \bArray_reg[5][18]  ( .D(n6221), .CK(clk), .RN(n7593), .Q(
        \bArray[5][18] ), .QN(n5416) );
  DFFRX1 \bArray_reg[3][18]  ( .D(n6317), .CK(clk), .RN(n7585), .Q(
        \bArray[3][18] ), .QN(n5512) );
  DFFRX1 \bArray_reg[7][18]  ( .D(n6125), .CK(clk), .RN(n7601), .Q(
        \bArray[7][18] ), .QN(n5320) );
  DFFRX1 \bArray_reg[0][18]  ( .D(n6461), .CK(clk), .RN(n7573), .Q(
        \bArray[0][18] ), .QN(n5656) );
  DFFRX1 \bArray_reg[4][18]  ( .D(n6269), .CK(clk), .RN(n7589), .Q(
        \bArray[4][18] ), .QN(n5464) );
  DFFRX1 \bArray_reg[2][17]  ( .D(n6364), .CK(clk), .RN(n7581), .Q(
        \bArray[2][17] ), .QN(n5559) );
  DFFRX1 \bArray_reg[6][17]  ( .D(n6172), .CK(clk), .RN(n7597), .Q(
        \bArray[6][17] ), .QN(n5367) );
  DFFRX1 \bArray_reg[10][18]  ( .D(n5981), .CK(clk), .RN(n7613), .Q(
        \bArray[10][18] ), .QN(n5176) );
  DFFRX1 \bArray_reg[10][17]  ( .D(n5980), .CK(clk), .RN(n7613), .Q(
        \bArray[10][17] ), .QN(n5175) );
  DFFRX1 \bArray_reg[14][18]  ( .D(n5789), .CK(clk), .RN(n7629), .Q(
        \bArray[14][18] ), .QN(n4984) );
  DFFRX1 \bArray_reg[14][17]  ( .D(n5788), .CK(clk), .RN(n7629), .Q(
        \bArray[14][17] ), .QN(n4983) );
  DFFRX1 \bArray_reg[1][17]  ( .D(n6412), .CK(clk), .RN(n7577), .Q(
        \bArray[1][17] ), .QN(n5607) );
  DFFRX1 \bArray_reg[5][17]  ( .D(n6220), .CK(clk), .RN(n7593), .Q(
        \bArray[5][17] ), .QN(n5415) );
  DFFRX1 \bArray_reg[9][18]  ( .D(n6029), .CK(clk), .RN(n7609), .Q(
        \bArray[9][18] ), .QN(n5224) );
  DFFRX1 \bArray_reg[9][17]  ( .D(n6028), .CK(clk), .RN(n7609), .Q(
        \bArray[9][17] ), .QN(n5223) );
  DFFRX1 \bArray_reg[13][18]  ( .D(n5837), .CK(clk), .RN(n7625), .Q(
        \bArray[13][18] ), .QN(n5032) );
  DFFRX1 \bArray_reg[13][17]  ( .D(n5836), .CK(clk), .RN(n7625), .Q(
        \bArray[13][17] ), .QN(n5031) );
  DFFRX1 \bArray_reg[3][17]  ( .D(n6316), .CK(clk), .RN(n7585), .Q(
        \bArray[3][17] ), .QN(n5511) );
  DFFRX1 \bArray_reg[7][17]  ( .D(n6124), .CK(clk), .RN(n7601), .Q(
        \bArray[7][17] ), .QN(n5319) );
  DFFRX1 \bArray_reg[11][18]  ( .D(n5933), .CK(clk), .RN(n7617), .Q(
        \bArray[11][18] ), .QN(n5128) );
  DFFRX1 \bArray_reg[11][17]  ( .D(n5932), .CK(clk), .RN(n7617), .Q(
        \bArray[11][17] ), .QN(n5127) );
  DFFRX1 \bArray_reg[15][18]  ( .D(n5741), .CK(clk), .RN(n7633), .Q(
        \bArray[15][18] ), .QN(n4936) );
  DFFRX1 \bArray_reg[15][17]  ( .D(n5740), .CK(clk), .RN(n7633), .Q(
        \bArray[15][17] ), .QN(n4935) );
  DFFRX1 \bArray_reg[0][17]  ( .D(n6460), .CK(clk), .RN(n7573), .Q(
        \bArray[0][17] ), .QN(n5655) );
  DFFRX1 \bArray_reg[4][17]  ( .D(n6268), .CK(clk), .RN(n7589), .Q(
        \bArray[4][17] ), .QN(n5463) );
  DFFRX1 \bArray_reg[8][18]  ( .D(n6077), .CK(clk), .RN(n7605), .Q(
        \bArray[8][18] ), .QN(n5272) );
  DFFRX1 \bArray_reg[8][17]  ( .D(n6076), .CK(clk), .RN(n7605), .Q(
        \bArray[8][17] ), .QN(n5271) );
  DFFRX1 \bArray_reg[12][18]  ( .D(n5885), .CK(clk), .RN(n7621), .Q(
        \bArray[12][18] ), .QN(n5080) );
  DFFRX1 \bArray_reg[12][17]  ( .D(n5884), .CK(clk), .RN(n7621), .Q(
        \bArray[12][17] ), .QN(n5079) );
  DFFRX1 \bArray_reg[2][16]  ( .D(n6363), .CK(clk), .RN(n7581), .Q(
        \bArray[2][16] ), .QN(n5558) );
  DFFRX1 \bArray_reg[10][16]  ( .D(n5979), .CK(clk), .RN(n7613), .Q(
        \bArray[10][16] ), .QN(n5174) );
  DFFRX1 \bArray_reg[1][16]  ( .D(n6411), .CK(clk), .RN(n7577), .Q(
        \bArray[1][16] ), .QN(n5606) );
  DFFRX1 \bArray_reg[5][16]  ( .D(n6219), .CK(clk), .RN(n7593), .Q(
        \bArray[5][16] ), .QN(n5414) );
  DFFRX1 \bArray_reg[9][16]  ( .D(n6027), .CK(clk), .RN(n7609), .Q(
        \bArray[9][16] ), .QN(n5222) );
  DFFRX1 \bArray_reg[13][16]  ( .D(n5835), .CK(clk), .RN(n7625), .Q(
        \bArray[13][16] ), .QN(n5030) );
  DFFRX1 \bArray_reg[3][16]  ( .D(n6315), .CK(clk), .RN(n7585), .Q(
        \bArray[3][16] ), .QN(n5510) );
  DFFRX1 \bArray_reg[11][16]  ( .D(n5931), .CK(clk), .RN(n7617), .Q(
        \bArray[11][16] ), .QN(n5126) );
  DFFRX1 \bArray_reg[0][16]  ( .D(n6459), .CK(clk), .RN(n7573), .Q(
        \bArray[0][16] ), .QN(n5654) );
  DFFRX1 \bArray_reg[4][16]  ( .D(n6267), .CK(clk), .RN(n7589), .Q(
        \bArray[4][16] ), .QN(n5462) );
  DFFRX1 \bArray_reg[8][16]  ( .D(n6075), .CK(clk), .RN(n7605), .Q(
        \bArray[8][16] ), .QN(n5270) );
  DFFRX1 \bArray_reg[12][16]  ( .D(n5883), .CK(clk), .RN(n7621), .Q(
        \bArray[12][16] ), .QN(n5078) );
  DFFRX1 \bArray_reg[6][16]  ( .D(n6171), .CK(clk), .RN(n7597), .Q(
        \bArray[6][16] ), .QN(n5366) );
  DFFRX1 \bArray_reg[14][16]  ( .D(n5787), .CK(clk), .RN(n7629), .Q(
        \bArray[14][16] ), .QN(n4982) );
  DFFRX1 \bArray_reg[7][16]  ( .D(n6123), .CK(clk), .RN(n7601), .Q(
        \bArray[7][16] ), .QN(n5318) );
  DFFRX1 \bArray_reg[15][16]  ( .D(n5739), .CK(clk), .RN(n7633), .Q(
        \bArray[15][16] ), .QN(n4934) );
  DFFQX1 \xArray_reg[8][9]  ( .D(N28266), .CK(clk), .Q(\xArray[8][9] ) );
  DFFQX1 \xArray_reg[2][9]  ( .D(N28650), .CK(clk), .Q(\xArray[2][9] ) );
  DFFQX1 \xArray_reg[8][8]  ( .D(N28265), .CK(clk), .Q(\xArray[8][8] ) );
  DFFQX1 \xArray_reg[8][7]  ( .D(N28264), .CK(clk), .Q(\xArray[8][7] ) );
  DFFQX1 \xArray_reg[2][8]  ( .D(N28649), .CK(clk), .Q(\xArray[2][8] ) );
  DFFQX1 \xArray_reg[2][7]  ( .D(N28648), .CK(clk), .Q(\xArray[2][7] ) );
  DFFQX1 \xArray_reg[8][6]  ( .D(N28263), .CK(clk), .Q(\xArray[8][6] ) );
  DFFQX1 \xArray_reg[8][5]  ( .D(N28262), .CK(clk), .Q(\xArray[8][5] ) );
  DFFQX1 \xArray_reg[2][6]  ( .D(N28647), .CK(clk), .Q(\xArray[2][6] ) );
  DFFQX1 \xArray_reg[8][1]  ( .D(N28258), .CK(clk), .Q(\xArray[8][1] ) );
  DFFQX1 \xArray_reg[8][0]  ( .D(N28257), .CK(clk), .Q(\xArray[8][0] ) );
  DFFQX1 \xArray_reg[8][2]  ( .D(N28259), .CK(clk), .Q(\xArray[8][2] ) );
  DFFQX1 \xArray_reg[8][3]  ( .D(N28260), .CK(clk), .Q(\xArray[8][3] ) );
  DFFQX1 \xArray_reg[2][5]  ( .D(N28646), .CK(clk), .Q(\xArray[2][5] ) );
  DFFQX1 \xArray_reg[2][4]  ( .D(N28645), .CK(clk), .Q(\xArray[2][4] ) );
  DFFQX1 \xArray_reg[2][1]  ( .D(N28642), .CK(clk), .Q(\xArray[2][1] ) );
  DFFQX1 \xArray_reg[2][3]  ( .D(N28644), .CK(clk), .Q(\xArray[2][3] ) );
  DFFQX1 \xArray_reg[2][0]  ( .D(N28641), .CK(clk), .Q(\xArray[2][0] ) );
  DFFQX1 \xArray_reg[14][55]  ( .D(N27928), .CK(clk), .Q(\xArray[14][55] ) );
  DFFQX1 \xArray_reg[10][55]  ( .D(N28184), .CK(clk), .Q(\xArray[10][55] ) );
  DFFQX1 \xArray_reg[10][54]  ( .D(N28183), .CK(clk), .Q(\xArray[10][54] ) );
  DFFQX1 \xArray_reg[6][55]  ( .D(N28440), .CK(clk), .Q(\xArray[6][55] ) );
  DFFQX1 \xArray_reg[6][54]  ( .D(N28439), .CK(clk), .Q(\xArray[6][54] ) );
  DFFQX1 \xArray_reg[14][54]  ( .D(N27927), .CK(clk), .Q(\xArray[14][54] ) );
  DFFQX1 \xArray_reg[14][53]  ( .D(N27926), .CK(clk), .Q(\xArray[14][53] ) );
  DFFQX1 \xArray_reg[14][52]  ( .D(N27925), .CK(clk), .Q(\xArray[14][52] ) );
  DFFQX1 \xArray_reg[10][53]  ( .D(N28182), .CK(clk), .Q(\xArray[10][53] ) );
  DFFQX1 \xArray_reg[10][52]  ( .D(N28181), .CK(clk), .Q(\xArray[10][52] ) );
  DFFQX1 \xArray_reg[6][53]  ( .D(N28438), .CK(clk), .Q(\xArray[6][53] ) );
  DFFQX1 \xArray_reg[6][52]  ( .D(N28437), .CK(clk), .Q(\xArray[6][52] ) );
  DFFQX1 \xArray_reg[14][51]  ( .D(N27924), .CK(clk), .Q(\xArray[14][51] ) );
  DFFQX1 \xArray_reg[10][51]  ( .D(N28180), .CK(clk), .Q(\xArray[10][51] ) );
  DFFQX1 \xArray_reg[10][50]  ( .D(N28179), .CK(clk), .Q(\xArray[10][50] ) );
  DFFQX1 \xArray_reg[6][51]  ( .D(N28436), .CK(clk), .Q(\xArray[6][51] ) );
  DFFQX1 \xArray_reg[6][50]  ( .D(N28435), .CK(clk), .Q(\xArray[6][50] ) );
  DFFQX1 \xArray_reg[14][50]  ( .D(N27923), .CK(clk), .Q(\xArray[14][50] ) );
  DFFQX1 \xArray_reg[10][49]  ( .D(N28178), .CK(clk), .Q(\xArray[10][49] ) );
  DFFQX1 \xArray_reg[6][49]  ( .D(N28434), .CK(clk), .Q(\xArray[6][49] ) );
  DFFQX1 \xArray_reg[3][34]  ( .D(N28611), .CK(clk), .Q(\xArray[3][34] ) );
  DFFQX1 \xArray_reg[4][33]  ( .D(N28546), .CK(clk), .Q(\xArray[4][33] ) );
  DFFQX1 \xArray_reg[15][9]  ( .D(N27818), .CK(clk), .Q(\xArray[15][9] ) );
  DFFQX1 \xArray_reg[14][9]  ( .D(N27882), .CK(clk), .Q(\xArray[14][9] ) );
  DFFQX1 \xArray_reg[5][9]  ( .D(N28458), .CK(clk), .Q(\xArray[5][9] ) );
  DFFQX1 \xArray_reg[5][8]  ( .D(N28457), .CK(clk), .Q(\xArray[5][8] ) );
  DFFQX1 \xArray_reg[4][9]  ( .D(N28522), .CK(clk), .Q(\xArray[4][9] ) );
  DFFQX1 \xArray_reg[11][8]  ( .D(N28073), .CK(clk), .Q(\xArray[11][8] ) );
  DFFQX1 \xArray_reg[12][8]  ( .D(N28009), .CK(clk), .Q(\xArray[12][8] ) );
  DFFQX1 \xArray_reg[7][8]  ( .D(N28329), .CK(clk), .Q(\xArray[7][8] ) );
  DFFQX1 \xArray_reg[10][8]  ( .D(N28137), .CK(clk), .Q(\xArray[10][8] ) );
  DFFQX1 \xArray_reg[6][8]  ( .D(N28393), .CK(clk), .Q(\xArray[6][8] ) );
  DFFQX1 \xArray_reg[9][9]  ( .D(N28202), .CK(clk), .Q(\xArray[9][9] ) );
  DFFQX1 \xArray_reg[3][9]  ( .D(N28586), .CK(clk), .Q(\xArray[3][9] ) );
  DFFQX1 \xArray_reg[3][8]  ( .D(N28585), .CK(clk), .Q(\xArray[3][8] ) );
  DFFQX1 \xArray_reg[14][8]  ( .D(N27881), .CK(clk), .Q(\xArray[14][8] ) );
  DFFQX1 \xArray_reg[14][7]  ( .D(N27880), .CK(clk), .Q(\xArray[14][7] ) );
  DFFQX1 \xArray_reg[0][8]  ( .D(N28777), .CK(clk), .Q(\xArray[0][8] ) );
  DFFQX1 \xArray_reg[5][7]  ( .D(N28456), .CK(clk), .Q(\xArray[5][7] ) );
  DFFQX1 \xArray_reg[4][7]  ( .D(N28520), .CK(clk), .Q(\xArray[4][7] ) );
  DFFQX1 \xArray_reg[4][8]  ( .D(N28521), .CK(clk), .Q(\xArray[4][8] ) );
  DFFQX1 \xArray_reg[11][7]  ( .D(N28072), .CK(clk), .Q(\xArray[11][7] ) );
  DFFQX1 \xArray_reg[12][7]  ( .D(N28008), .CK(clk), .Q(\xArray[12][7] ) );
  DFFQX1 \xArray_reg[11][6]  ( .D(N28071), .CK(clk), .Q(\xArray[11][6] ) );
  DFFQX1 \xArray_reg[12][6]  ( .D(N28007), .CK(clk), .Q(\xArray[12][6] ) );
  DFFQX1 \xArray_reg[7][6]  ( .D(N28327), .CK(clk), .Q(\xArray[7][6] ) );
  DFFQX1 \xArray_reg[1][8]  ( .D(N28713), .CK(clk), .Q(\xArray[1][8] ) );
  DFFQX1 \xArray_reg[1][7]  ( .D(N28712), .CK(clk), .Q(\xArray[1][7] ) );
  DFFQX1 \xArray_reg[13][8]  ( .D(N27945), .CK(clk), .Q(\xArray[13][8] ) );
  DFFQX1 \xArray_reg[13][7]  ( .D(N27944), .CK(clk), .Q(\xArray[13][7] ) );
  DFFQX1 \xArray_reg[9][8]  ( .D(N28201), .CK(clk), .Q(\xArray[9][8] ) );
  DFFQX1 \xArray_reg[3][6]  ( .D(N28583), .CK(clk), .Q(\xArray[3][6] ) );
  DFFQX1 \xArray_reg[15][5]  ( .D(N27814), .CK(clk), .Q(\xArray[15][5] ) );
  DFFQX1 \xArray_reg[0][5]  ( .D(N28774), .CK(clk), .Q(\xArray[0][5] ) );
  DFFQX1 \xArray_reg[14][6]  ( .D(N27879), .CK(clk), .Q(\xArray[14][6] ) );
  DFFQX1 \xArray_reg[14][5]  ( .D(N27878), .CK(clk), .Q(\xArray[14][5] ) );
  DFFQX1 \xArray_reg[5][5]  ( .D(N28454), .CK(clk), .Q(\xArray[5][5] ) );
  DFFQX1 \xArray_reg[4][6]  ( .D(N28519), .CK(clk), .Q(\xArray[4][6] ) );
  DFFQX1 \xArray_reg[4][5]  ( .D(N28518), .CK(clk), .Q(\xArray[4][5] ) );
  DFFQX1 \xArray_reg[11][5]  ( .D(N28070), .CK(clk), .Q(\xArray[11][5] ) );
  DFFQX1 \xArray_reg[11][4]  ( .D(N28069), .CK(clk), .Q(\xArray[11][4] ) );
  DFFQX1 \xArray_reg[11][3]  ( .D(N28068), .CK(clk), .Q(\xArray[11][3] ) );
  DFFQX1 \xArray_reg[12][5]  ( .D(N28006), .CK(clk), .Q(\xArray[12][5] ) );
  DFFQX1 \xArray_reg[12][4]  ( .D(N28005), .CK(clk), .Q(\xArray[12][4] ) );
  DFFQX1 \xArray_reg[12][3]  ( .D(N28004), .CK(clk), .Q(\xArray[12][3] ) );
  DFFQX1 \xArray_reg[7][5]  ( .D(N28326), .CK(clk), .Q(\xArray[7][5] ) );
  DFFQX1 \xArray_reg[1][6]  ( .D(N28711), .CK(clk), .Q(\xArray[1][6] ) );
  DFFQX1 \xArray_reg[1][5]  ( .D(N28710), .CK(clk), .Q(\xArray[1][5] ) );
  DFFQX1 \xArray_reg[13][6]  ( .D(N27943), .CK(clk), .Q(\xArray[13][6] ) );
  DFFQX1 \xArray_reg[13][5]  ( .D(N27942), .CK(clk), .Q(\xArray[13][5] ) );
  DFFQX1 \xArray_reg[10][6]  ( .D(N28135), .CK(clk), .Q(\xArray[10][6] ) );
  DFFQX1 \xArray_reg[10][5]  ( .D(N28134), .CK(clk), .Q(\xArray[10][5] ) );
  DFFQX1 \xArray_reg[6][6]  ( .D(N28391), .CK(clk), .Q(\xArray[6][6] ) );
  DFFQX1 \xArray_reg[6][5]  ( .D(N28390), .CK(clk), .Q(\xArray[6][5] ) );
  DFFQX1 \xArray_reg[9][5]  ( .D(N28198), .CK(clk), .Q(\xArray[9][5] ) );
  DFFQX1 \xArray_reg[3][5]  ( .D(N28582), .CK(clk), .Q(\xArray[3][5] ) );
  DFFQX1 \xArray_reg[3][4]  ( .D(N28581), .CK(clk), .Q(\xArray[3][4] ) );
  DFFQX1 \xArray_reg[3][2]  ( .D(N28579), .CK(clk), .Q(\xArray[3][2] ) );
  DFFQX1 \xArray_reg[3][0]  ( .D(N28577), .CK(clk), .Q(\xArray[3][0] ) );
  DFFQX1 \xArray_reg[3][3]  ( .D(N28580), .CK(clk), .Q(\xArray[3][3] ) );
  DFFQX1 \xArray_reg[15][4]  ( .D(N27813), .CK(clk), .Q(\xArray[15][4] ) );
  DFFQX1 \xArray_reg[15][3]  ( .D(N27812), .CK(clk), .Q(\xArray[15][3] ) );
  DFFQX1 \xArray_reg[15][2]  ( .D(N27811), .CK(clk), .Q(\xArray[15][2] ) );
  DFFQX1 \xArray_reg[15][1]  ( .D(N27810), .CK(clk), .Q(\xArray[15][1] ) );
  DFFQX1 \xArray_reg[15][0]  ( .D(N27809), .CK(clk), .Q(\xArray[15][0] ) );
  DFFQX1 \xArray_reg[14][1]  ( .D(N27874), .CK(clk), .Q(\xArray[14][1] ) );
  DFFQX1 \xArray_reg[14][0]  ( .D(N27873), .CK(clk), .Q(\xArray[14][0] ) );
  DFFQX1 \xArray_reg[0][4]  ( .D(N28773), .CK(clk), .Q(\xArray[0][4] ) );
  DFFQX1 \xArray_reg[0][3]  ( .D(N28772), .CK(clk), .Q(\xArray[0][3] ) );
  DFFQX1 \xArray_reg[0][1]  ( .D(N28770), .CK(clk), .Q(\xArray[0][1] ) );
  DFFQX1 \xArray_reg[0][2]  ( .D(N28771), .CK(clk), .Q(\xArray[0][2] ) );
  DFFQX1 \xArray_reg[0][0]  ( .D(N28769), .CK(clk), .Q(\xArray[0][0] ) );
  DFFQX1 \xArray_reg[14][3]  ( .D(N27876), .CK(clk), .Q(\xArray[14][3] ) );
  DFFQX1 \xArray_reg[3][1]  ( .D(N28578), .CK(clk), .Q(\xArray[3][1] ) );
  DFFQX1 \xArray_reg[5][4]  ( .D(N28453), .CK(clk), .Q(\xArray[5][4] ) );
  DFFQX1 \xArray_reg[5][3]  ( .D(N28452), .CK(clk), .Q(\xArray[5][3] ) );
  DFFQX1 \xArray_reg[5][1]  ( .D(N28450), .CK(clk), .Q(\xArray[5][1] ) );
  DFFQX1 \xArray_reg[5][0]  ( .D(N28449), .CK(clk), .Q(\xArray[5][0] ) );
  DFFQX1 \xArray_reg[4][4]  ( .D(N28517), .CK(clk), .Q(\xArray[4][4] ) );
  DFFQX1 \xArray_reg[4][2]  ( .D(N28515), .CK(clk), .Q(\xArray[4][2] ) );
  DFFQX1 \xArray_reg[4][1]  ( .D(N28514), .CK(clk), .Q(\xArray[4][1] ) );
  DFFQX1 \xArray_reg[4][0]  ( .D(N28513), .CK(clk), .Q(\xArray[4][0] ) );
  DFFQX1 \xArray_reg[11][0]  ( .D(N28065), .CK(clk), .Q(\xArray[11][0] ) );
  DFFQX1 \xArray_reg[11][1]  ( .D(N28066), .CK(clk), .Q(\xArray[11][1] ) );
  DFFQX1 \xArray_reg[12][1]  ( .D(N28002), .CK(clk), .Q(\xArray[12][1] ) );
  DFFQX1 \xArray_reg[12][0]  ( .D(N28001), .CK(clk), .Q(\xArray[12][0] ) );
  DFFQX1 \xArray_reg[7][0]  ( .D(N28321), .CK(clk), .Q(\xArray[7][0] ) );
  DFFQX1 \xArray_reg[7][4]  ( .D(N28325), .CK(clk), .Q(\xArray[7][4] ) );
  DFFQX1 \xArray_reg[7][3]  ( .D(N28324), .CK(clk), .Q(\xArray[7][3] ) );
  DFFQX1 \xArray_reg[7][2]  ( .D(N28323), .CK(clk), .Q(\xArray[7][2] ) );
  DFFQX1 \xArray_reg[7][1]  ( .D(N28322), .CK(clk), .Q(\xArray[7][1] ) );
  DFFQX1 \xArray_reg[14][2]  ( .D(N27875), .CK(clk), .Q(\xArray[14][2] ) );
  DFFQX1 \xArray_reg[12][2]  ( .D(N28003), .CK(clk), .Q(\xArray[12][2] ) );
  DFFQX1 \xArray_reg[5][2]  ( .D(N28451), .CK(clk), .Q(\xArray[5][2] ) );
  DFFQX1 \xArray_reg[1][4]  ( .D(N28709), .CK(clk), .Q(\xArray[1][4] ) );
  DFFQX1 \xArray_reg[1][1]  ( .D(N28706), .CK(clk), .Q(\xArray[1][1] ) );
  DFFQX1 \xArray_reg[1][3]  ( .D(N28708), .CK(clk), .Q(\xArray[1][3] ) );
  DFFQX1 \xArray_reg[1][0]  ( .D(N28705), .CK(clk), .Q(\xArray[1][0] ) );
  DFFQX1 \xArray_reg[13][4]  ( .D(N27941), .CK(clk), .Q(\xArray[13][4] ) );
  DFFQX1 \xArray_reg[13][3]  ( .D(N27940), .CK(clk), .Q(\xArray[13][3] ) );
  DFFQX1 \xArray_reg[13][0]  ( .D(N27937), .CK(clk), .Q(\xArray[13][0] ) );
  DFFQX1 \xArray_reg[10][1]  ( .D(N28130), .CK(clk), .Q(\xArray[10][1] ) );
  DFFQX1 \xArray_reg[10][0]  ( .D(N28129), .CK(clk), .Q(\xArray[10][0] ) );
  DFFQX1 \xArray_reg[10][4]  ( .D(N28133), .CK(clk), .Q(\xArray[10][4] ) );
  DFFQX1 \xArray_reg[6][0]  ( .D(N28385), .CK(clk), .Q(\xArray[6][0] ) );
  DFFQX1 \xArray_reg[6][4]  ( .D(N28389), .CK(clk), .Q(\xArray[6][4] ) );
  DFFQX1 \xArray_reg[6][3]  ( .D(N28388), .CK(clk), .Q(\xArray[6][3] ) );
  DFFQX1 \xArray_reg[6][1]  ( .D(N28386), .CK(clk), .Q(\xArray[6][1] ) );
  DFFQX1 \xArray_reg[9][4]  ( .D(N28197), .CK(clk), .Q(\xArray[9][4] ) );
  DFFQX1 \xArray_reg[9][3]  ( .D(N28196), .CK(clk), .Q(\xArray[9][3] ) );
  DFFQX1 \xArray_reg[9][1]  ( .D(N28194), .CK(clk), .Q(\xArray[9][1] ) );
  DFFQX1 \xArray_reg[9][0]  ( .D(N28193), .CK(clk), .Q(\xArray[9][0] ) );
  DFFQX1 \xArray_reg[1][2]  ( .D(N28707), .CK(clk), .Q(\xArray[1][2] ) );
  DFFQX1 \xArray_reg[10][2]  ( .D(N28131), .CK(clk), .Q(\xArray[10][2] ) );
  DFFQX1 \xArray_reg[13][2]  ( .D(N27939), .CK(clk), .Q(\xArray[13][2] ) );
  DFFQX1 \xArray_reg[9][2]  ( .D(N28195), .CK(clk), .Q(\xArray[9][2] ) );
  DFFRX4 \xCount_reg[3]  ( .D(xCount_next[3]), .CK(clk), .RN(n7639), .Q(N1764), 
        .QN(n106) );
  DFFQX1 \xArray_reg[9][26]  ( .D(N28219), .CK(clk), .Q(\xArray[9][26] ) );
  DFFQX1 \xArray_reg[9][24]  ( .D(N28217), .CK(clk), .Q(\xArray[9][24] ) );
  DFFQX1 \xArray_reg[9][25]  ( .D(N28218), .CK(clk), .Q(\xArray[9][25] ) );
  DFFQX1 \xArray_reg[6][24]  ( .D(N28409), .CK(clk), .Q(\xArray[6][24] ) );
  DFFQX1 \xArray_reg[8][24]  ( .D(N28281), .CK(clk), .Q(\xArray[8][24] ) );
  DFFQX1 \xArray_reg[2][26]  ( .D(N28667), .CK(clk), .Q(\xArray[2][26] ) );
  DFFQX1 \xArray_reg[2][25]  ( .D(N28666), .CK(clk), .Q(\xArray[2][25] ) );
  DFFQX1 \xArray_reg[3][26]  ( .D(N28603), .CK(clk), .Q(\xArray[3][26] ) );
  DFFQX1 \xArray_reg[14][26]  ( .D(N27899), .CK(clk), .Q(\xArray[14][26] ) );
  DFFQX1 \xArray_reg[14][25]  ( .D(N27898), .CK(clk), .Q(\xArray[14][25] ) );
  DFFQX1 \xArray_reg[1][23]  ( .D(N28728), .CK(clk), .Q(\xArray[1][23] ) );
  DFFQX1 \xArray_reg[13][23]  ( .D(N27960), .CK(clk), .Q(\xArray[13][23] ) );
  DFFQX1 \xArray_reg[10][23]  ( .D(N28152), .CK(clk), .Q(\xArray[10][23] ) );
  DFFQX1 \xArray_reg[10][22]  ( .D(N28151), .CK(clk), .Q(\xArray[10][22] ) );
  DFFQX1 \xArray_reg[1][24]  ( .D(N28729), .CK(clk), .Q(\xArray[1][24] ) );
  DFFQX1 \xArray_reg[6][22]  ( .D(N28407), .CK(clk), .Q(\xArray[6][22] ) );
  DFFQX1 \xArray_reg[13][24]  ( .D(N27961), .CK(clk), .Q(\xArray[13][24] ) );
  DFFQX1 \xArray_reg[9][23]  ( .D(N28216), .CK(clk), .Q(\xArray[9][23] ) );
  DFFQX1 \xArray_reg[9][22]  ( .D(N28215), .CK(clk), .Q(\xArray[9][22] ) );
  DFFQX1 \xArray_reg[6][23]  ( .D(N28408), .CK(clk), .Q(\xArray[6][23] ) );
  DFFQX1 \xArray_reg[8][23]  ( .D(N28280), .CK(clk), .Q(\xArray[8][23] ) );
  DFFQX1 \xArray_reg[8][22]  ( .D(N28279), .CK(clk), .Q(\xArray[8][22] ) );
  DFFQX1 \xArray_reg[2][23]  ( .D(N28664), .CK(clk), .Q(\xArray[2][23] ) );
  DFFQX1 \xArray_reg[2][24]  ( .D(N28665), .CK(clk), .Q(\xArray[2][24] ) );
  DFFQX1 \xArray_reg[3][25]  ( .D(N28602), .CK(clk), .Q(\xArray[3][25] ) );
  DFFQX1 \xArray_reg[15][23]  ( .D(N27832), .CK(clk), .Q(\xArray[15][23] ) );
  DFFQX1 \xArray_reg[14][23]  ( .D(N27896), .CK(clk), .Q(\xArray[14][23] ) );
  DFFQX1 \xArray_reg[14][24]  ( .D(N27897), .CK(clk), .Q(\xArray[14][24] ) );
  DFFQX1 \xArray_reg[0][23]  ( .D(N28792), .CK(clk), .Q(\xArray[0][23] ) );
  DFFQX1 \xArray_reg[5][23]  ( .D(N28472), .CK(clk), .Q(\xArray[5][23] ) );
  DFFQX1 \xArray_reg[4][23]  ( .D(N28536), .CK(clk), .Q(\xArray[4][23] ) );
  DFFQX1 \xArray_reg[11][22]  ( .D(N28087), .CK(clk), .Q(\xArray[11][22] ) );
  DFFQX1 \xArray_reg[11][23]  ( .D(N28088), .CK(clk), .Q(\xArray[11][23] ) );
  DFFQX1 \xArray_reg[12][23]  ( .D(N28024), .CK(clk), .Q(\xArray[12][23] ) );
  DFFQX1 \xArray_reg[12][22]  ( .D(N28023), .CK(clk), .Q(\xArray[12][22] ) );
  DFFQX1 \xArray_reg[7][22]  ( .D(N28343), .CK(clk), .Q(\xArray[7][22] ) );
  DFFQX1 \xArray_reg[7][23]  ( .D(N28344), .CK(clk), .Q(\xArray[7][23] ) );
  DFFQX1 \xArray_reg[1][22]  ( .D(N28727), .CK(clk), .Q(\xArray[1][22] ) );
  DFFQX1 \xArray_reg[13][22]  ( .D(N27959), .CK(clk), .Q(\xArray[13][22] ) );
  DFFQX1 \xArray_reg[10][21]  ( .D(N28150), .CK(clk), .Q(\xArray[10][21] ) );
  DFFQX1 \xArray_reg[6][21]  ( .D(N28406), .CK(clk), .Q(\xArray[6][21] ) );
  DFFQX1 \xArray_reg[9][21]  ( .D(N28214), .CK(clk), .Q(\xArray[9][21] ) );
  DFFQX1 \xArray_reg[8][21]  ( .D(N28278), .CK(clk), .Q(\xArray[8][21] ) );
  DFFQX1 \xArray_reg[2][22]  ( .D(N28663), .CK(clk), .Q(\xArray[2][22] ) );
  DFFQX1 \xArray_reg[3][23]  ( .D(N28600), .CK(clk), .Q(\xArray[3][23] ) );
  DFFQX1 \xArray_reg[15][22]  ( .D(N27831), .CK(clk), .Q(\xArray[15][22] ) );
  DFFQX1 \xArray_reg[14][22]  ( .D(N27895), .CK(clk), .Q(\xArray[14][22] ) );
  DFFQX1 \xArray_reg[0][22]  ( .D(N28791), .CK(clk), .Q(\xArray[0][22] ) );
  DFFQX1 \xArray_reg[5][22]  ( .D(N28471), .CK(clk), .Q(\xArray[5][22] ) );
  DFFQX1 \xArray_reg[5][21]  ( .D(N28470), .CK(clk), .Q(\xArray[5][21] ) );
  DFFQX1 \xArray_reg[4][22]  ( .D(N28535), .CK(clk), .Q(\xArray[4][22] ) );
  DFFQX1 \xArray_reg[11][21]  ( .D(N28086), .CK(clk), .Q(\xArray[11][21] ) );
  DFFQX1 \xArray_reg[12][21]  ( .D(N28022), .CK(clk), .Q(\xArray[12][21] ) );
  DFFQX1 \xArray_reg[7][21]  ( .D(N28342), .CK(clk), .Q(\xArray[7][21] ) );
  DFFQXL \xArray_reg[15][32]  ( .D(N27841), .CK(clk), .Q(\xArray[15][32] ) );
  DFFQXL \xArray_reg[0][32]  ( .D(N28801), .CK(clk), .Q(\xArray[0][32] ) );
  DFFQXL \xArray_reg[4][32]  ( .D(N28545), .CK(clk), .Q(\xArray[4][32] ) );
  DFFQXL \xArray_reg[11][32]  ( .D(N28097), .CK(clk), .Q(\xArray[11][32] ) );
  DFFQXL \xArray_reg[12][32]  ( .D(N28033), .CK(clk), .Q(\xArray[12][32] ) );
  DFFQXL \xArray_reg[7][32]  ( .D(N28353), .CK(clk), .Q(\xArray[7][32] ) );
  DFFQX1 \xArray_reg[2][30]  ( .D(N28671), .CK(clk), .Q(\xArray[2][30] ) );
  DFFQX1 \xArray_reg[2][29]  ( .D(N28670), .CK(clk), .Q(\xArray[2][29] ) );
  DFFQX1 \xArray_reg[2][63]  ( .D(N28704), .CK(clk), .Q(\xArray[2][63] ) );
  DFFQX1 \xArray_reg[2][62]  ( .D(N28703), .CK(clk), .Q(\xArray[2][62] ) );
  DFFQX1 \xArray_reg[2][61]  ( .D(N28702), .CK(clk), .Q(\xArray[2][61] ) );
  DFFQX1 \xArray_reg[2][60]  ( .D(N28701), .CK(clk), .Q(\xArray[2][60] ) );
  DFFQX1 \xArray_reg[2][59]  ( .D(N28700), .CK(clk), .Q(\xArray[2][59] ) );
  DFFQX1 \xArray_reg[2][58]  ( .D(N28699), .CK(clk), .Q(\xArray[2][58] ) );
  DFFQX1 \xArray_reg[2][57]  ( .D(N28698), .CK(clk), .Q(\xArray[2][57] ) );
  DFFQX1 \xArray_reg[2][56]  ( .D(N28697), .CK(clk), .Q(\xArray[2][56] ) );
  DFFQX1 \xArray_reg[14][63]  ( .D(N27936), .CK(clk), .Q(\xArray[14][63] ) );
  DFFQX1 \xArray_reg[10][63]  ( .D(N28192), .CK(clk), .Q(\xArray[10][63] ) );
  DFFQX1 \xArray_reg[6][63]  ( .D(N28448), .CK(clk), .Q(\xArray[6][63] ) );
  DFFQX1 \xArray_reg[10][62]  ( .D(N28191), .CK(clk), .Q(\xArray[10][62] ) );
  DFFQX1 \xArray_reg[6][62]  ( .D(N28447), .CK(clk), .Q(\xArray[6][62] ) );
  DFFQX1 \xArray_reg[14][62]  ( .D(N27935), .CK(clk), .Q(\xArray[14][62] ) );
  DFFQX1 \xArray_reg[14][61]  ( .D(N27934), .CK(clk), .Q(\xArray[14][61] ) );
  DFFQX1 \xArray_reg[10][61]  ( .D(N28190), .CK(clk), .Q(\xArray[10][61] ) );
  DFFQX1 \xArray_reg[6][61]  ( .D(N28446), .CK(clk), .Q(\xArray[6][61] ) );
  DFFQX1 \xArray_reg[14][60]  ( .D(N27933), .CK(clk), .Q(\xArray[14][60] ) );
  DFFQX1 \xArray_reg[10][59]  ( .D(N28188), .CK(clk), .Q(\xArray[10][59] ) );
  DFFQX1 \xArray_reg[10][60]  ( .D(N28189), .CK(clk), .Q(\xArray[10][60] ) );
  DFFQX1 \xArray_reg[6][60]  ( .D(N28445), .CK(clk), .Q(\xArray[6][60] ) );
  DFFQX1 \xArray_reg[6][59]  ( .D(N28444), .CK(clk), .Q(\xArray[6][59] ) );
  DFFQX1 \xArray_reg[14][59]  ( .D(N27932), .CK(clk), .Q(\xArray[14][59] ) );
  DFFQX1 \xArray_reg[14][58]  ( .D(N27931), .CK(clk), .Q(\xArray[14][58] ) );
  DFFQX1 \xArray_reg[10][58]  ( .D(N28187), .CK(clk), .Q(\xArray[10][58] ) );
  DFFQX1 \xArray_reg[6][58]  ( .D(N28443), .CK(clk), .Q(\xArray[6][58] ) );
  DFFQX1 \xArray_reg[14][57]  ( .D(N27930), .CK(clk), .Q(\xArray[14][57] ) );
  DFFQX1 \xArray_reg[10][57]  ( .D(N28186), .CK(clk), .Q(\xArray[10][57] ) );
  DFFQX1 \xArray_reg[10][56]  ( .D(N28185), .CK(clk), .Q(\xArray[10][56] ) );
  DFFQX1 \xArray_reg[6][57]  ( .D(N28442), .CK(clk), .Q(\xArray[6][57] ) );
  DFFQX1 \xArray_reg[6][56]  ( .D(N28441), .CK(clk), .Q(\xArray[6][56] ) );
  DFFQX1 \xArray_reg[14][56]  ( .D(N27929), .CK(clk), .Q(\xArray[14][56] ) );
  DFFRX1 out_valid_reg ( .D(N35192), .CK(clk), .RN(n7647), .QN(n6689) );
  DFFRX1 \x_out_reg[0]  ( .D(N34942), .CK(clk), .RN(n7644), .QN(n6687) );
  DFFRX1 \x_out_reg[1]  ( .D(N34943), .CK(clk), .RN(n7644), .QN(n6685) );
  DFFRX1 \x_out_reg[2]  ( .D(N34944), .CK(clk), .RN(n7644), .QN(n6683) );
  DFFRX1 \x_out_reg[3]  ( .D(N34945), .CK(clk), .RN(n7644), .QN(n6681) );
  DFFRX1 \x_out_reg[4]  ( .D(N34946), .CK(clk), .RN(n7644), .QN(n6679) );
  DFFRX1 \x_out_reg[5]  ( .D(N34947), .CK(clk), .RN(n7644), .QN(n6677) );
  DFFRX1 \x_out_reg[6]  ( .D(N34948), .CK(clk), .RN(n7644), .QN(n6675) );
  DFFRX1 \x_out_reg[7]  ( .D(N34949), .CK(clk), .RN(n7644), .QN(n6673) );
  DFFRX1 \x_out_reg[8]  ( .D(N34950), .CK(clk), .RN(n7644), .QN(n6671) );
  DFFRX1 \x_out_reg[9]  ( .D(N34951), .CK(clk), .RN(n7644), .QN(n6669) );
  DFFRX1 \x_out_reg[10]  ( .D(N34952), .CK(clk), .RN(n7644), .QN(n6667) );
  DFFRX1 \x_out_reg[11]  ( .D(N34953), .CK(clk), .RN(n7643), .QN(n6665) );
  DFFRX1 \x_out_reg[12]  ( .D(N34954), .CK(clk), .RN(n7643), .QN(n6663) );
  DFFRX1 \x_out_reg[13]  ( .D(N34955), .CK(clk), .RN(n7643), .QN(n6661) );
  DFFRX1 \x_out_reg[14]  ( .D(N34956), .CK(clk), .RN(n7643), .QN(n6659) );
  DFFRX1 \x_out_reg[15]  ( .D(N34957), .CK(clk), .RN(n7643), .QN(n6657) );
  DFFRX1 \x_out_reg[16]  ( .D(N34958), .CK(clk), .RN(n7643), .QN(n6655) );
  DFFRX1 \x_out_reg[17]  ( .D(N34959), .CK(clk), .RN(n7643), .QN(n6653) );
  DFFRX1 \x_out_reg[18]  ( .D(N34960), .CK(clk), .RN(n7643), .QN(n6651) );
  DFFRX1 \x_out_reg[19]  ( .D(N34961), .CK(clk), .RN(n7643), .QN(n6649) );
  DFFRX1 \x_out_reg[20]  ( .D(N34962), .CK(clk), .RN(n7643), .QN(n6647) );
  DFFRX1 \x_out_reg[21]  ( .D(N34963), .CK(clk), .RN(n7643), .QN(n6645) );
  DFFRX1 \x_out_reg[22]  ( .D(N34964), .CK(clk), .RN(n7643), .QN(n6643) );
  DFFRX1 \x_out_reg[23]  ( .D(N34965), .CK(clk), .RN(n7642), .QN(n6641) );
  DFFRX1 \x_out_reg[24]  ( .D(N34966), .CK(clk), .RN(n7642), .QN(n6639) );
  DFFRX1 \x_out_reg[25]  ( .D(N34967), .CK(clk), .RN(n7642), .QN(n6637) );
  DFFRX1 \x_out_reg[26]  ( .D(N34968), .CK(clk), .RN(n7642), .QN(n6635) );
  DFFRX1 \x_out_reg[27]  ( .D(N34969), .CK(clk), .RN(n7642), .QN(n6633) );
  DFFRX1 \x_out_reg[28]  ( .D(N34970), .CK(clk), .RN(n7642), .QN(n6631) );
  DFFRX1 \x_out_reg[29]  ( .D(N34971), .CK(clk), .RN(n7642), .QN(n6629) );
  DFFRX1 \x_out_reg[30]  ( .D(N34972), .CK(clk), .RN(n7642), .QN(n6627) );
  DFFRX1 \x_out_reg[31]  ( .D(N34973), .CK(clk), .RN(n7642), .QN(n6625) );
  DFFQX1 \xArray_reg[8][4]  ( .D(N28261), .CK(clk), .Q(\xArray[8][4] ) );
  DFFQX1 \xArray_reg[3][7]  ( .D(N28584), .CK(clk), .Q(\xArray[3][7] ) );
  DFFQX1 \xArray_reg[7][7]  ( .D(N28328), .CK(clk), .Q(\xArray[7][7] ) );
  DFFQX1 \xArray_reg[9][7]  ( .D(N28200), .CK(clk), .Q(\xArray[9][7] ) );
  DFFQX1 \xArray_reg[10][7]  ( .D(N28136), .CK(clk), .Q(\xArray[10][7] ) );
  DFFQX1 \xArray_reg[6][7]  ( .D(N28392), .CK(clk), .Q(\xArray[6][7] ) );
  DFFQX1 \xArray_reg[15][7]  ( .D(N27816), .CK(clk), .Q(\xArray[15][7] ) );
  DFFQX1 \xArray_reg[0][7]  ( .D(N28776), .CK(clk), .Q(\xArray[0][7] ) );
  DFFQX1 \xArray_reg[4][3]  ( .D(N28516), .CK(clk), .Q(\xArray[4][3] ) );
  DFFQX1 \xArray_reg[10][3]  ( .D(N28132), .CK(clk), .Q(\xArray[10][3] ) );
  DFFQX1 \xArray_reg[0][9]  ( .D(N28778), .CK(clk), .Q(\xArray[0][9] ) );
  DFFQX1 \xArray_reg[11][9]  ( .D(N28074), .CK(clk), .Q(\xArray[11][9] ) );
  DFFQX1 \xArray_reg[12][9]  ( .D(N28010), .CK(clk), .Q(\xArray[12][9] ) );
  DFFQX1 \xArray_reg[7][9]  ( .D(N28330), .CK(clk), .Q(\xArray[7][9] ) );
  DFFQX1 \xArray_reg[1][9]  ( .D(N28714), .CK(clk), .Q(\xArray[1][9] ) );
  DFFQX1 \xArray_reg[13][9]  ( .D(N27946), .CK(clk), .Q(\xArray[13][9] ) );
  DFFQX1 \xArray_reg[10][9]  ( .D(N28138), .CK(clk), .Q(\xArray[10][9] ) );
  DFFQX1 \xArray_reg[6][9]  ( .D(N28394), .CK(clk), .Q(\xArray[6][9] ) );
  DFFQX1 \xArray_reg[15][6]  ( .D(N27815), .CK(clk), .Q(\xArray[15][6] ) );
  DFFQX1 \xArray_reg[0][6]  ( .D(N28775), .CK(clk), .Q(\xArray[0][6] ) );
  DFFQX1 \xArray_reg[14][4]  ( .D(N27877), .CK(clk), .Q(\xArray[14][4] ) );
  DFFQX1 \xArray_reg[13][1]  ( .D(N27938), .CK(clk), .Q(\xArray[13][1] ) );
  DFFQX1 \xArray_reg[8][20]  ( .D(N28277), .CK(clk), .Q(\xArray[8][20] ) );
  DFFQX1 \xArray_reg[3][22]  ( .D(N28599), .CK(clk), .Q(\xArray[3][22] ) );
  DFFQX1 \xArray_reg[15][21]  ( .D(N27830), .CK(clk), .Q(\xArray[15][21] ) );
  DFFQX1 \xArray_reg[14][21]  ( .D(N27894), .CK(clk), .Q(\xArray[14][21] ) );
  DFFQX1 \xArray_reg[0][21]  ( .D(N28790), .CK(clk), .Q(\xArray[0][21] ) );
  DFFQX1 \xArray_reg[4][21]  ( .D(N28534), .CK(clk), .Q(\xArray[4][21] ) );
  DFFQX1 \xArray_reg[12][20]  ( .D(N28021), .CK(clk), .Q(\xArray[12][20] ) );
  DFFQX1 \xArray_reg[13][21]  ( .D(N27958), .CK(clk), .Q(\xArray[13][21] ) );
  DFFQX1 \xArray_reg[10][20]  ( .D(N28149), .CK(clk), .Q(\xArray[10][20] ) );
  DFFQX1 \xArray_reg[6][20]  ( .D(N28405), .CK(clk), .Q(\xArray[6][20] ) );
  DFFQX1 \xArray_reg[9][20]  ( .D(N28213), .CK(clk), .Q(\xArray[9][20] ) );
  DFFQX1 \xArray_reg[1][20]  ( .D(N28725), .CK(clk), .Q(\xArray[1][20] ) );
  DFFQX1 \xArray_reg[1][21]  ( .D(N28726), .CK(clk), .Q(\xArray[1][21] ) );
  DFFQX1 \xArray_reg[1][19]  ( .D(N28724), .CK(clk), .Q(\xArray[1][19] ) );
  DFFQX1 \xArray_reg[13][20]  ( .D(N27957), .CK(clk), .Q(\xArray[13][20] ) );
  DFFQX1 \xArray_reg[13][19]  ( .D(N27956), .CK(clk), .Q(\xArray[13][19] ) );
  DFFQX1 \xArray_reg[10][19]  ( .D(N28148), .CK(clk), .Q(\xArray[10][19] ) );
  DFFQX1 \xArray_reg[10][18]  ( .D(N28147), .CK(clk), .Q(\xArray[10][18] ) );
  DFFQX1 \xArray_reg[6][19]  ( .D(N28404), .CK(clk), .Q(\xArray[6][19] ) );
  DFFQX1 \xArray_reg[6][18]  ( .D(N28403), .CK(clk), .Q(\xArray[6][18] ) );
  DFFQX1 \xArray_reg[9][19]  ( .D(N28212), .CK(clk), .Q(\xArray[9][19] ) );
  DFFQX1 \xArray_reg[8][19]  ( .D(N28276), .CK(clk), .Q(\xArray[8][19] ) );
  DFFQX1 \xArray_reg[8][18]  ( .D(N28275), .CK(clk), .Q(\xArray[8][18] ) );
  DFFQX1 \xArray_reg[2][20]  ( .D(N28661), .CK(clk), .Q(\xArray[2][20] ) );
  DFFQX1 \xArray_reg[2][19]  ( .D(N28660), .CK(clk), .Q(\xArray[2][19] ) );
  DFFQX1 \xArray_reg[2][21]  ( .D(N28662), .CK(clk), .Q(\xArray[2][21] ) );
  DFFQX1 \xArray_reg[3][21]  ( .D(N28598), .CK(clk), .Q(\xArray[3][21] ) );
  DFFQX1 \xArray_reg[3][20]  ( .D(N28597), .CK(clk), .Q(\xArray[3][20] ) );
  DFFQX1 \xArray_reg[15][19]  ( .D(N27828), .CK(clk), .Q(\xArray[15][19] ) );
  DFFQX1 \xArray_reg[15][20]  ( .D(N27829), .CK(clk), .Q(\xArray[15][20] ) );
  DFFQX1 \xArray_reg[14][20]  ( .D(N27893), .CK(clk), .Q(\xArray[14][20] ) );
  DFFQX1 \xArray_reg[14][19]  ( .D(N27892), .CK(clk), .Q(\xArray[14][19] ) );
  DFFQX1 \xArray_reg[0][20]  ( .D(N28789), .CK(clk), .Q(\xArray[0][20] ) );
  DFFQX1 \xArray_reg[0][19]  ( .D(N28788), .CK(clk), .Q(\xArray[0][19] ) );
  DFFQX1 \xArray_reg[5][20]  ( .D(N28469), .CK(clk), .Q(\xArray[5][20] ) );
  DFFQX1 \xArray_reg[5][19]  ( .D(N28468), .CK(clk), .Q(\xArray[5][19] ) );
  DFFQX1 \xArray_reg[4][20]  ( .D(N28533), .CK(clk), .Q(\xArray[4][20] ) );
  DFFQX1 \xArray_reg[4][19]  ( .D(N28532), .CK(clk), .Q(\xArray[4][19] ) );
  DFFQX1 \xArray_reg[11][19]  ( .D(N28084), .CK(clk), .Q(\xArray[11][19] ) );
  DFFQX1 \xArray_reg[11][20]  ( .D(N28085), .CK(clk), .Q(\xArray[11][20] ) );
  DFFQX1 \xArray_reg[12][19]  ( .D(N28020), .CK(clk), .Q(\xArray[12][19] ) );
  DFFQX1 \xArray_reg[7][19]  ( .D(N28340), .CK(clk), .Q(\xArray[7][19] ) );
  DFFQX1 \xArray_reg[7][20]  ( .D(N28341), .CK(clk), .Q(\xArray[7][20] ) );
  DFFQX1 \xArray_reg[1][17]  ( .D(N28722), .CK(clk), .Q(\xArray[1][17] ) );
  DFFQX1 \xArray_reg[1][18]  ( .D(N28723), .CK(clk), .Q(\xArray[1][18] ) );
  DFFQX1 \xArray_reg[13][17]  ( .D(N27954), .CK(clk), .Q(\xArray[13][17] ) );
  DFFQX1 \xArray_reg[13][18]  ( .D(N27955), .CK(clk), .Q(\xArray[13][18] ) );
  DFFQX1 \xArray_reg[10][17]  ( .D(N28146), .CK(clk), .Q(\xArray[10][17] ) );
  DFFQX1 \xArray_reg[6][17]  ( .D(N28402), .CK(clk), .Q(\xArray[6][17] ) );
  DFFQX1 \xArray_reg[9][18]  ( .D(N28211), .CK(clk), .Q(\xArray[9][18] ) );
  DFFQX1 \xArray_reg[9][17]  ( .D(N28210), .CK(clk), .Q(\xArray[9][17] ) );
  DFFQX1 \xArray_reg[8][17]  ( .D(N28274), .CK(clk), .Q(\xArray[8][17] ) );
  DFFQX1 \xArray_reg[8][16]  ( .D(N28273), .CK(clk), .Q(\xArray[8][16] ) );
  DFFQX1 \xArray_reg[2][17]  ( .D(N28658), .CK(clk), .Q(\xArray[2][17] ) );
  DFFQX1 \xArray_reg[2][18]  ( .D(N28659), .CK(clk), .Q(\xArray[2][18] ) );
  DFFQX1 \xArray_reg[3][19]  ( .D(N28596), .CK(clk), .Q(\xArray[3][19] ) );
  DFFQX1 \xArray_reg[3][18]  ( .D(N28595), .CK(clk), .Q(\xArray[3][18] ) );
  DFFQX1 \xArray_reg[15][18]  ( .D(N27827), .CK(clk), .Q(\xArray[15][18] ) );
  DFFQX1 \xArray_reg[15][17]  ( .D(N27826), .CK(clk), .Q(\xArray[15][17] ) );
  DFFQX1 \xArray_reg[14][18]  ( .D(N27891), .CK(clk), .Q(\xArray[14][18] ) );
  DFFQX1 \xArray_reg[0][18]  ( .D(N28787), .CK(clk), .Q(\xArray[0][18] ) );
  DFFQX1 \xArray_reg[0][17]  ( .D(N28786), .CK(clk), .Q(\xArray[0][17] ) );
  DFFQX1 \xArray_reg[5][18]  ( .D(N28467), .CK(clk), .Q(\xArray[5][18] ) );
  DFFQX1 \xArray_reg[5][17]  ( .D(N28466), .CK(clk), .Q(\xArray[5][17] ) );
  DFFQX1 \xArray_reg[4][18]  ( .D(N28531), .CK(clk), .Q(\xArray[4][18] ) );
  DFFQX1 \xArray_reg[4][17]  ( .D(N28530), .CK(clk), .Q(\xArray[4][17] ) );
  DFFQX1 \xArray_reg[11][17]  ( .D(N28082), .CK(clk), .Q(\xArray[11][17] ) );
  DFFQX1 \xArray_reg[11][18]  ( .D(N28083), .CK(clk), .Q(\xArray[11][18] ) );
  DFFQX1 \xArray_reg[12][17]  ( .D(N28018), .CK(clk), .Q(\xArray[12][17] ) );
  DFFQX1 \xArray_reg[12][18]  ( .D(N28019), .CK(clk), .Q(\xArray[12][18] ) );
  DFFQX1 \xArray_reg[7][17]  ( .D(N28338), .CK(clk), .Q(\xArray[7][17] ) );
  DFFQX1 \xArray_reg[7][18]  ( .D(N28339), .CK(clk), .Q(\xArray[7][18] ) );
  DFFQX1 \xArray_reg[1][16]  ( .D(N28721), .CK(clk), .Q(\xArray[1][16] ) );
  DFFQX1 \xArray_reg[13][16]  ( .D(N27953), .CK(clk), .Q(\xArray[13][16] ) );
  DFFQX1 \xArray_reg[10][16]  ( .D(N28145), .CK(clk), .Q(\xArray[10][16] ) );
  DFFQX1 \xArray_reg[10][15]  ( .D(N28144), .CK(clk), .Q(\xArray[10][15] ) );
  DFFQX1 \xArray_reg[6][16]  ( .D(N28401), .CK(clk), .Q(\xArray[6][16] ) );
  DFFQX1 \xArray_reg[6][15]  ( .D(N28400), .CK(clk), .Q(\xArray[6][15] ) );
  DFFQX1 \xArray_reg[9][16]  ( .D(N28209), .CK(clk), .Q(\xArray[9][16] ) );
  DFFQX1 \xArray_reg[9][15]  ( .D(N28208), .CK(clk), .Q(\xArray[9][15] ) );
  DFFQX1 \xArray_reg[8][15]  ( .D(N28272), .CK(clk), .Q(\xArray[8][15] ) );
  DFFQX1 \xArray_reg[2][16]  ( .D(N28657), .CK(clk), .Q(\xArray[2][16] ) );
  DFFQX1 \xArray_reg[2][15]  ( .D(N28656), .CK(clk), .Q(\xArray[2][15] ) );
  DFFQX1 \xArray_reg[3][16]  ( .D(N28593), .CK(clk), .Q(\xArray[3][16] ) );
  DFFQX1 \xArray_reg[3][17]  ( .D(N28594), .CK(clk), .Q(\xArray[3][17] ) );
  DFFQX1 \xArray_reg[15][15]  ( .D(N27824), .CK(clk), .Q(\xArray[15][15] ) );
  DFFQX1 \xArray_reg[15][16]  ( .D(N27825), .CK(clk), .Q(\xArray[15][16] ) );
  DFFQX1 \xArray_reg[14][16]  ( .D(N27889), .CK(clk), .Q(\xArray[14][16] ) );
  DFFQX1 \xArray_reg[14][17]  ( .D(N27890), .CK(clk), .Q(\xArray[14][17] ) );
  DFFQX1 \xArray_reg[5][15]  ( .D(N28464), .CK(clk), .Q(\xArray[5][15] ) );
  DFFQX1 \xArray_reg[5][16]  ( .D(N28465), .CK(clk), .Q(\xArray[5][16] ) );
  DFFQX1 \xArray_reg[4][16]  ( .D(N28529), .CK(clk), .Q(\xArray[4][16] ) );
  DFFQX1 \xArray_reg[11][15]  ( .D(N28080), .CK(clk), .Q(\xArray[11][15] ) );
  DFFQX1 \xArray_reg[12][16]  ( .D(N28017), .CK(clk), .Q(\xArray[12][16] ) );
  DFFQX1 \xArray_reg[12][15]  ( .D(N28016), .CK(clk), .Q(\xArray[12][15] ) );
  DFFQX1 \xArray_reg[11][16]  ( .D(N28081), .CK(clk), .Q(\xArray[11][16] ) );
  DFFQX1 \xArray_reg[7][16]  ( .D(N28337), .CK(clk), .Q(\xArray[7][16] ) );
  DFFQX1 \xArray_reg[7][15]  ( .D(N28336), .CK(clk), .Q(\xArray[7][15] ) );
  DFFQX1 \xArray_reg[8][13]  ( .D(N28270), .CK(clk), .Q(\xArray[8][13] ) );
  DFFQX1 \xArray_reg[8][14]  ( .D(N28271), .CK(clk), .Q(\xArray[8][14] ) );
  DFFQX1 \xArray_reg[2][14]  ( .D(N28655), .CK(clk), .Q(\xArray[2][14] ) );
  DFFQX1 \xArray_reg[3][15]  ( .D(N28592), .CK(clk), .Q(\xArray[3][15] ) );
  DFFQX1 \xArray_reg[3][14]  ( .D(N28591), .CK(clk), .Q(\xArray[3][14] ) );
  DFFQX1 \xArray_reg[15][13]  ( .D(N27822), .CK(clk), .Q(\xArray[15][13] ) );
  DFFQX1 \xArray_reg[15][14]  ( .D(N27823), .CK(clk), .Q(\xArray[15][14] ) );
  DFFQX1 \xArray_reg[14][14]  ( .D(N27887), .CK(clk), .Q(\xArray[14][14] ) );
  DFFQX1 \xArray_reg[14][15]  ( .D(N27888), .CK(clk), .Q(\xArray[14][15] ) );
  DFFQX1 \xArray_reg[5][13]  ( .D(N28462), .CK(clk), .Q(\xArray[5][13] ) );
  DFFQX1 \xArray_reg[5][14]  ( .D(N28463), .CK(clk), .Q(\xArray[5][14] ) );
  DFFQX1 \xArray_reg[4][14]  ( .D(N28527), .CK(clk), .Q(\xArray[4][14] ) );
  DFFQX1 \xArray_reg[4][15]  ( .D(N28528), .CK(clk), .Q(\xArray[4][15] ) );
  DFFQX1 \xArray_reg[11][13]  ( .D(N28078), .CK(clk), .Q(\xArray[11][13] ) );
  DFFQX1 \xArray_reg[11][14]  ( .D(N28079), .CK(clk), .Q(\xArray[11][14] ) );
  DFFQX1 \xArray_reg[12][13]  ( .D(N28014), .CK(clk), .Q(\xArray[12][13] ) );
  DFFQX1 \xArray_reg[12][14]  ( .D(N28015), .CK(clk), .Q(\xArray[12][14] ) );
  DFFQX1 \xArray_reg[7][13]  ( .D(N28334), .CK(clk), .Q(\xArray[7][13] ) );
  DFFQX1 \xArray_reg[7][14]  ( .D(N28335), .CK(clk), .Q(\xArray[7][14] ) );
  DFFQX1 \xArray_reg[1][14]  ( .D(N28719), .CK(clk), .Q(\xArray[1][14] ) );
  DFFQX1 \xArray_reg[1][15]  ( .D(N28720), .CK(clk), .Q(\xArray[1][15] ) );
  DFFQX1 \xArray_reg[13][14]  ( .D(N27951), .CK(clk), .Q(\xArray[13][14] ) );
  DFFQX1 \xArray_reg[13][15]  ( .D(N27952), .CK(clk), .Q(\xArray[13][15] ) );
  DFFQX1 \xArray_reg[10][13]  ( .D(N28142), .CK(clk), .Q(\xArray[10][13] ) );
  DFFQX1 \xArray_reg[10][14]  ( .D(N28143), .CK(clk), .Q(\xArray[10][14] ) );
  DFFQX1 \xArray_reg[6][13]  ( .D(N28398), .CK(clk), .Q(\xArray[6][13] ) );
  DFFQX1 \xArray_reg[6][14]  ( .D(N28399), .CK(clk), .Q(\xArray[6][14] ) );
  DFFQX1 \xArray_reg[9][13]  ( .D(N28206), .CK(clk), .Q(\xArray[9][13] ) );
  DFFQX1 \xArray_reg[9][14]  ( .D(N28207), .CK(clk), .Q(\xArray[9][14] ) );
  DFFQX1 \xArray_reg[8][11]  ( .D(N28268), .CK(clk), .Q(\xArray[8][11] ) );
  DFFQX1 \xArray_reg[8][12]  ( .D(N28269), .CK(clk), .Q(\xArray[8][12] ) );
  DFFQX1 \xArray_reg[2][12]  ( .D(N28653), .CK(clk), .Q(\xArray[2][12] ) );
  DFFQX1 \xArray_reg[2][13]  ( .D(N28654), .CK(clk), .Q(\xArray[2][13] ) );
  DFFQX1 \xArray_reg[3][12]  ( .D(N28589), .CK(clk), .Q(\xArray[3][12] ) );
  DFFQX1 \xArray_reg[3][13]  ( .D(N28590), .CK(clk), .Q(\xArray[3][13] ) );
  DFFQX1 \xArray_reg[15][12]  ( .D(N27821), .CK(clk), .Q(\xArray[15][12] ) );
  DFFQX1 \xArray_reg[14][12]  ( .D(N27885), .CK(clk), .Q(\xArray[14][12] ) );
  DFFQX1 \xArray_reg[14][13]  ( .D(N27886), .CK(clk), .Q(\xArray[14][13] ) );
  DFFQX1 \xArray_reg[5][12]  ( .D(N28461), .CK(clk), .Q(\xArray[5][12] ) );
  DFFQX1 \xArray_reg[5][11]  ( .D(N28460), .CK(clk), .Q(\xArray[5][11] ) );
  DFFQX1 \xArray_reg[4][13]  ( .D(N28526), .CK(clk), .Q(\xArray[4][13] ) );
  DFFQX1 \xArray_reg[4][12]  ( .D(N28525), .CK(clk), .Q(\xArray[4][12] ) );
  DFFQX1 \xArray_reg[11][12]  ( .D(N28077), .CK(clk), .Q(\xArray[11][12] ) );
  DFFQX1 \xArray_reg[12][12]  ( .D(N28013), .CK(clk), .Q(\xArray[12][12] ) );
  DFFQX1 \xArray_reg[11][11]  ( .D(N28076), .CK(clk), .Q(\xArray[11][11] ) );
  DFFQX1 \xArray_reg[12][11]  ( .D(N28012), .CK(clk), .Q(\xArray[12][11] ) );
  DFFQX1 \xArray_reg[7][11]  ( .D(N28332), .CK(clk), .Q(\xArray[7][11] ) );
  DFFQX1 \xArray_reg[7][12]  ( .D(N28333), .CK(clk), .Q(\xArray[7][12] ) );
  DFFQX1 \xArray_reg[1][13]  ( .D(N28718), .CK(clk), .Q(\xArray[1][13] ) );
  DFFQX1 \xArray_reg[1][12]  ( .D(N28717), .CK(clk), .Q(\xArray[1][12] ) );
  DFFQX1 \xArray_reg[13][13]  ( .D(N27950), .CK(clk), .Q(\xArray[13][13] ) );
  DFFQX1 \xArray_reg[13][12]  ( .D(N27949), .CK(clk), .Q(\xArray[13][12] ) );
  DFFQX1 \xArray_reg[10][12]  ( .D(N28141), .CK(clk), .Q(\xArray[10][12] ) );
  DFFQX1 \xArray_reg[10][11]  ( .D(N28140), .CK(clk), .Q(\xArray[10][11] ) );
  DFFQX1 \xArray_reg[6][12]  ( .D(N28397), .CK(clk), .Q(\xArray[6][12] ) );
  DFFQX1 \xArray_reg[6][11]  ( .D(N28396), .CK(clk), .Q(\xArray[6][11] ) );
  DFFQX1 \xArray_reg[9][12]  ( .D(N28205), .CK(clk), .Q(\xArray[9][12] ) );
  DFFQX1 \xArray_reg[9][11]  ( .D(N28204), .CK(clk), .Q(\xArray[9][11] ) );
  DFFQX1 \xArray_reg[8][10]  ( .D(N28267), .CK(clk), .Q(\xArray[8][10] ) );
  DFFQX1 \xArray_reg[2][11]  ( .D(N28652), .CK(clk), .Q(\xArray[2][11] ) );
  DFFQX1 \xArray_reg[2][10]  ( .D(N28651), .CK(clk), .Q(\xArray[2][10] ) );
  DFFQX1 \xArray_reg[3][11]  ( .D(N28588), .CK(clk), .Q(\xArray[3][11] ) );
  DFFQX1 \xArray_reg[15][10]  ( .D(N27819), .CK(clk), .Q(\xArray[15][10] ) );
  DFFQX1 \xArray_reg[15][11]  ( .D(N27820), .CK(clk), .Q(\xArray[15][11] ) );
  DFFQX1 \xArray_reg[14][11]  ( .D(N27884), .CK(clk), .Q(\xArray[14][11] ) );
  DFFQX1 \xArray_reg[14][10]  ( .D(N27883), .CK(clk), .Q(\xArray[14][10] ) );
  DFFQX1 \xArray_reg[0][11]  ( .D(N28780), .CK(clk), .Q(\xArray[0][11] ) );
  DFFQX1 \xArray_reg[0][10]  ( .D(N28779), .CK(clk), .Q(\xArray[0][10] ) );
  DFFQX1 \xArray_reg[5][10]  ( .D(N28459), .CK(clk), .Q(\xArray[5][10] ) );
  DFFQX1 \xArray_reg[4][11]  ( .D(N28524), .CK(clk), .Q(\xArray[4][11] ) );
  DFFQX1 \xArray_reg[4][10]  ( .D(N28523), .CK(clk), .Q(\xArray[4][10] ) );
  DFFQX1 \xArray_reg[11][10]  ( .D(N28075), .CK(clk), .Q(\xArray[11][10] ) );
  DFFQX1 \xArray_reg[12][10]  ( .D(N28011), .CK(clk), .Q(\xArray[12][10] ) );
  DFFQX1 \xArray_reg[7][10]  ( .D(N28331), .CK(clk), .Q(\xArray[7][10] ) );
  DFFQX1 \xArray_reg[1][11]  ( .D(N28716), .CK(clk), .Q(\xArray[1][11] ) );
  DFFQX1 \xArray_reg[1][10]  ( .D(N28715), .CK(clk), .Q(\xArray[1][10] ) );
  DFFQX1 \xArray_reg[13][11]  ( .D(N27948), .CK(clk), .Q(\xArray[13][11] ) );
  DFFQX1 \xArray_reg[13][10]  ( .D(N27947), .CK(clk), .Q(\xArray[13][10] ) );
  DFFQX1 \xArray_reg[10][10]  ( .D(N28139), .CK(clk), .Q(\xArray[10][10] ) );
  DFFQX1 \xArray_reg[6][10]  ( .D(N28395), .CK(clk), .Q(\xArray[6][10] ) );
  DFFQX1 \xArray_reg[9][10]  ( .D(N28203), .CK(clk), .Q(\xArray[9][10] ) );
  DFFQX1 \xArray_reg[3][10]  ( .D(N28587), .CK(clk), .Q(\xArray[3][10] ) );
  DFFQX1 \xArray_reg[11][2]  ( .D(N28067), .CK(clk), .Q(\xArray[11][2] ) );
  DFFQX1 \xArray_reg[6][2]  ( .D(N28387), .CK(clk), .Q(\xArray[6][2] ) );
  DFFQX1 \xArray_reg[2][2]  ( .D(N28643), .CK(clk), .Q(\xArray[2][2] ) );
  DFFQX1 \xArray_reg[3][33]  ( .D(N28610), .CK(clk), .Q(\xArray[3][33] ) );
  DFFQX1 \xArray_reg[3][32]  ( .D(N28609), .CK(clk), .Q(\xArray[3][32] ) );
  DFFQX1 \xArray_reg[3][31]  ( .D(N28608), .CK(clk), .Q(\xArray[3][31] ) );
  DFFQX1 \xArray_reg[3][30]  ( .D(N28607), .CK(clk), .Q(\xArray[3][30] ) );
  DFFQX1 \xArray_reg[3][29]  ( .D(N28606), .CK(clk), .Q(\xArray[3][29] ) );
  DFFQX1 \xArray_reg[2][28]  ( .D(N28669), .CK(clk), .Q(\xArray[2][28] ) );
  DFFQX1 \xArray_reg[2][27]  ( .D(N28668), .CK(clk), .Q(\xArray[2][27] ) );
  DFFQX1 \xArray_reg[5][32]  ( .D(N28481), .CK(clk), .Q(\xArray[5][32] ) );
  DFFQX1 \xArray_reg[14][29]  ( .D(N27902), .CK(clk), .Q(\xArray[14][29] ) );
  DFFQX1 \xArray_reg[14][28]  ( .D(N27901), .CK(clk), .Q(\xArray[14][28] ) );
  DFFQX1 \xArray_reg[3][28]  ( .D(N28605), .CK(clk), .Q(\xArray[3][28] ) );
  DFFQX1 \xArray_reg[3][27]  ( .D(N28604), .CK(clk), .Q(\xArray[3][27] ) );
  DFFQX1 \xArray_reg[14][27]  ( .D(N27900), .CK(clk), .Q(\xArray[14][27] ) );
  DFFQX1 \xArray_reg[9][27]  ( .D(N28220), .CK(clk), .Q(\xArray[9][27] ) );
  DFFQX1 \xArray_reg[9][6]  ( .D(N28199), .CK(clk), .Q(\xArray[9][6] ) );
  DFFQX1 \xArray_reg[5][6]  ( .D(N28455), .CK(clk), .Q(\xArray[5][6] ) );
  OA22XL U7371 ( .A0(n7760), .A1(n727), .B0(n8350), .B1(n1262), .Y(n1261) );
  OR3X6 U7372 ( .A(n6698), .B(n6699), .C(n6622), .Y(N33773) );
  OAI222XL U7373 ( .A0(n8080), .A1(n3027), .B0(n8018), .B1(n3379), .C0(n8068), 
        .C1(n3098), .Y(n3951) );
  OAI222XL U7374 ( .A0(n8080), .A1(n3026), .B0(n8018), .B1(n3378), .C0(n3149), 
        .C1(n3097), .Y(n3933) );
  INVX1 U7375 ( .A(n2543), .Y(n8515) );
  INVX1 U7376 ( .A(n2371), .Y(n8514) );
  OAI222XL U7377 ( .A0(n8083), .A1(n3023), .B0(n8019), .B1(n3375), .C0(n8070), 
        .C1(n3094), .Y(n3879) );
  INVX1 U7378 ( .A(n2540), .Y(n8500) );
  INVX1 U7379 ( .A(n2362), .Y(n8499) );
  OAI222XL U7380 ( .A0(n8083), .A1(n3022), .B0(n8019), .B1(n3374), .C0(n8070), 
        .C1(n3093), .Y(n3861) );
  INVX1 U7381 ( .A(n2539), .Y(n8495) );
  INVX1 U7382 ( .A(n2359), .Y(n8494) );
  OAI222X1 U7383 ( .A0(n8083), .A1(n3014), .B0(n8019), .B1(n3366), .C0(n8070), 
        .C1(n3085), .Y(n3717) );
  INVX3 U7384 ( .A(\xArray[14][3] ), .Y(n9374) );
  OA22X1 U7385 ( .A0(n7757), .A1(n638), .B0(n8346), .B1(n923), .Y(n922) );
  OAI221X1 U7386 ( .A0(\xArray[6][17] ), .A1(n8293), .B0(\xArray[10][17] ), 
        .B1(n8239), .C0(n1483), .Y(n923) );
  OA22X1 U7387 ( .A0(n7746), .A1(n558), .B0(n8346), .B1(n893), .Y(n892) );
  OA22X1 U7388 ( .A0(n7750), .A1(n478), .B0(n8337), .B1(n863), .Y(n862) );
  OA22X1 U7389 ( .A0(n7741), .A1(n398), .B0(n8345), .B1(n833), .Y(n832) );
  OA22X1 U7390 ( .A0(n7755), .A1(n1182), .B0(n8344), .B1(n1676), .Y(n1675) );
  OA22X1 U7391 ( .A0(n7759), .A1(n711), .B0(n8350), .B1(n1252), .Y(n1251) );
  OA22X1 U7392 ( .A0(n7759), .A1(n719), .B0(n8350), .B1(n1257), .Y(n1256) );
  NAND3X4 U7393 ( .A(n6696), .B(n6697), .C(n1266), .Y(N33903) );
  OA22X1 U7394 ( .A0(n7760), .A1(n735), .B0(n8350), .B1(n1267), .Y(n1266) );
  OA22X1 U7395 ( .A0(n7753), .A1(n950), .B0(n8341), .B1(n1518), .Y(n1517) );
  NAND3X1 U7396 ( .A(n6691), .B(n6692), .C(n1725), .Y(n1262) );
  OA22X1 U7397 ( .A0(n7753), .A1(n959), .B0(n8340), .B1(n1530), .Y(n1529) );
  OA22X1 U7398 ( .A0(n7745), .A1(n1132), .B0(n8344), .B1(n1646), .Y(n1645) );
  CLKBUFX3 U7399 ( .A(n7226), .Y(n7225) );
  OA22X1 U7400 ( .A0(n7745), .A1(n1082), .B0(n8343), .B1(n1616), .Y(n1615) );
  OA22X1 U7401 ( .A0(n7754), .A1(n1032), .B0(n8343), .B1(n1586), .Y(n1585) );
  MX4X1 U7402 ( .A(n7015), .B(n7013), .C(n7014), .D(n7012), .S0(n7224), .S1(
        n7223), .Y(N28879) );
  MX4X1 U7403 ( .A(n7019), .B(n7017), .C(n7018), .D(n7016), .S0(n7224), .S1(
        n7223), .Y(N28878) );
  MX4X1 U7404 ( .A(n7023), .B(n7021), .C(n7022), .D(n7020), .S0(n7224), .S1(
        n7223), .Y(N28877) );
  MX4X1 U7405 ( .A(n7027), .B(n7025), .C(n7026), .D(n7024), .S0(n7224), .S1(
        n7223), .Y(N28876) );
  MX4X1 U7406 ( .A(n7031), .B(n7029), .C(n7030), .D(n7028), .S0(n7224), .S1(
        n7223), .Y(N28875) );
  MX4X1 U7407 ( .A(\bArray[0][21] ), .B(\bArray[1][21] ), .C(\bArray[2][21] ), 
        .D(\bArray[3][21] ), .S0(n7207), .S1(n7219), .Y(n7031) );
  MX4X1 U7408 ( .A(n7047), .B(n7045), .C(n7046), .D(n7044), .S0(n7225), .S1(
        n7223), .Y(N28871) );
  MX4X1 U7409 ( .A(n7043), .B(n7041), .C(n7042), .D(n7040), .S0(n7224), .S1(
        n7223), .Y(N28872) );
  MX4X1 U7410 ( .A(n7039), .B(n7037), .C(n7038), .D(n7036), .S0(n7224), .S1(
        n7223), .Y(N28873) );
  MX4X1 U7411 ( .A(n7035), .B(n7033), .C(n7034), .D(n7032), .S0(n7224), .S1(
        n7223), .Y(N28874) );
  NAND3X4 U7412 ( .A(n6701), .B(n6702), .C(n1271), .Y(N33902) );
  OAI221X1 U7413 ( .A0(\xArray[5][3] ), .A1(n8280), .B0(\xArray[9][3] ), .B1(
        n8226), .C0(n1734), .Y(n1277) );
  CLKBUFX3 U7414 ( .A(n7739), .Y(n7715) );
  CLKBUFX3 U7415 ( .A(n8219), .Y(n8204) );
  OA22X1 U7416 ( .A0(n7755), .A1(n1232), .B0(n8345), .B1(n1706), .Y(n1705) );
  MX4X1 U7417 ( .A(n7051), .B(n7049), .C(n7050), .D(n7048), .S0(n7225), .S1(
        n8408), .Y(N28870) );
  MX4X1 U7418 ( .A(n7055), .B(n7053), .C(n7054), .D(n7052), .S0(n7225), .S1(
        n8408), .Y(N28869) );
  MX4X1 U7419 ( .A(n7059), .B(n7057), .C(n7058), .D(n7056), .S0(n7225), .S1(
        n8408), .Y(N28868) );
  MX4X1 U7420 ( .A(n7063), .B(n7061), .C(n7062), .D(n7060), .S0(n7225), .S1(
        n8408), .Y(N28867) );
  MX4X1 U7421 ( .A(n7067), .B(n7065), .C(n7066), .D(n7064), .S0(n7225), .S1(
        n8408), .Y(N28866) );
  MX4X1 U7422 ( .A(n7071), .B(n7069), .C(n7070), .D(n7068), .S0(n7225), .S1(
        n8408), .Y(N28865) );
  MX4X1 U7423 ( .A(n7075), .B(n7073), .C(n7074), .D(n7072), .S0(n7225), .S1(
        n8408), .Y(N28864) );
  MX4X1 U7424 ( .A(n7083), .B(n7081), .C(n7082), .D(n7080), .S0(n7225), .S1(
        n8408), .Y(N28862) );
  MX4X1 U7425 ( .A(n7079), .B(n7077), .C(n7078), .D(n7076), .S0(n7225), .S1(
        n8408), .Y(N28863) );
  MX4X1 U7426 ( .A(n7087), .B(n7085), .C(n7086), .D(n7084), .S0(n7225), .S1(
        n8885), .Y(N28861) );
  MX4X1 U7427 ( .A(n7091), .B(n7089), .C(n7090), .D(n7088), .S0(n7225), .S1(
        n8885), .Y(N28860) );
  MX4X1 U7428 ( .A(n7095), .B(n7093), .C(n7094), .D(n7092), .S0(n7225), .S1(
        n8885), .Y(N28859) );
  MX4X1 U7429 ( .A(n7099), .B(n7097), .C(n7098), .D(n7096), .S0(n8407), .S1(
        N1763), .Y(N28858) );
  MX4X1 U7430 ( .A(n7103), .B(n7101), .C(n7102), .D(n7100), .S0(n8407), .S1(
        N1763), .Y(N28857) );
  MX4X1 U7431 ( .A(n7107), .B(n7105), .C(n7106), .D(n7104), .S0(n8407), .S1(
        N1763), .Y(N28856) );
  MX4X1 U7432 ( .A(n7111), .B(n7109), .C(n7110), .D(n7108), .S0(n8407), .S1(
        N1763), .Y(N28855) );
  MX4X1 U7433 ( .A(n7115), .B(n7113), .C(n7114), .D(n7112), .S0(n8407), .S1(
        N1763), .Y(N28854) );
  MX4X1 U7434 ( .A(n7119), .B(n7117), .C(n7118), .D(n7116), .S0(n7226), .S1(
        N1763), .Y(N28853) );
  MX4X1 U7435 ( .A(n7123), .B(n7121), .C(n7122), .D(n7120), .S0(n7226), .S1(
        N1763), .Y(N28852) );
  MX4X1 U7436 ( .A(n7127), .B(n7125), .C(n7126), .D(n7124), .S0(n7226), .S1(
        N1763), .Y(N28851) );
  MX4X1 U7437 ( .A(n7131), .B(n7129), .C(n7130), .D(n7128), .S0(n7226), .S1(
        N1763), .Y(N28850) );
  MX4X1 U7438 ( .A(n7135), .B(n7133), .C(n7134), .D(n7132), .S0(n7226), .S1(
        n7223), .Y(N28849) );
  MX4X1 U7439 ( .A(n7139), .B(n7137), .C(n7138), .D(n7136), .S0(n7224), .S1(
        n8408), .Y(N28848) );
  MX4X1 U7440 ( .A(n7143), .B(n7141), .C(n7142), .D(n7140), .S0(n6700), .S1(
        n8408), .Y(N28847) );
  MX4X1 U7441 ( .A(n7151), .B(n7149), .C(n7150), .D(n7148), .S0(n7227), .S1(
        n8408), .Y(N28845) );
  MX4X1 U7442 ( .A(n7147), .B(n7145), .C(n7146), .D(n7144), .S0(n6700), .S1(
        n8408), .Y(N28846) );
  MX4X1 U7443 ( .A(n7155), .B(n7153), .C(n7154), .D(n7152), .S0(n7227), .S1(
        n8885), .Y(N28844) );
  MX4X1 U7444 ( .A(n7159), .B(n7157), .C(n7158), .D(n7156), .S0(n7227), .S1(
        n8885), .Y(N28843) );
  MX4X1 U7445 ( .A(n7163), .B(n7161), .C(n7162), .D(n7160), .S0(n7227), .S1(
        n8885), .Y(N28842) );
  MX4X1 U7446 ( .A(n7167), .B(n7165), .C(n7166), .D(n7164), .S0(n7227), .S1(
        N1763), .Y(N28841) );
  MX4X1 U7447 ( .A(n7171), .B(n7169), .C(n7170), .D(n7168), .S0(n7227), .S1(
        N1763), .Y(N28840) );
  OAI221X1 U7448 ( .A0(\xArray[7][23] ), .A1(n8297), .B0(\xArray[11][23] ), 
        .B1(n8243), .C0(n1179), .Y(n589) );
  OAI221X1 U7449 ( .A0(\xArray[5][2] ), .A1(n8280), .B0(\xArray[9][2] ), .B1(
        n8226), .C0(n1737), .Y(n1282) );
  OAI211X1 U7450 ( .A0(n7742), .A1(n1492), .B0(n2189), .C0(n2190), .Y(N33720)
         );
  NAND2BX1 U7451 ( .AN(n656), .B(n657), .Y(N34040) );
  OAI211X1 U7452 ( .A0(n7747), .A1(n1484), .B0(n2171), .C0(n2172), .Y(N33722)
         );
  OAI211X1 U7453 ( .A0(n7747), .A1(n1488), .B0(n2180), .C0(n2181), .Y(N33721)
         );
  NAND2BX1 U7454 ( .AN(n640), .B(n641), .Y(N34042) );
  NAND2BX1 U7455 ( .AN(n648), .B(n649), .Y(N34041) );
  OAI211X1 U7456 ( .A0(n7747), .A1(n1480), .B0(n2162), .C0(n2163), .Y(N33723)
         );
  NAND2BX1 U7457 ( .AN(n632), .B(n633), .Y(N34043) );
  OAI211X1 U7458 ( .A0(n7747), .A1(n1476), .B0(n2153), .C0(n2154), .Y(N33724)
         );
  NAND2BX1 U7459 ( .AN(n624), .B(n625), .Y(N34044) );
  OAI211X1 U7460 ( .A0(n7745), .A1(n1472), .B0(n2144), .C0(n2145), .Y(N33725)
         );
  NAND2BX1 U7461 ( .AN(n616), .B(n617), .Y(N34045) );
  OAI211X1 U7462 ( .A0(n7747), .A1(n1468), .B0(n2135), .C0(n2136), .Y(N33726)
         );
  NAND2BX1 U7463 ( .AN(n608), .B(n609), .Y(N34046) );
  OAI211X1 U7464 ( .A0(n7743), .A1(n1464), .B0(n2126), .C0(n2127), .Y(N33727)
         );
  NAND2BX1 U7465 ( .AN(n600), .B(n601), .Y(N34047) );
  OAI211X1 U7466 ( .A0(n7743), .A1(n1448), .B0(n2090), .C0(n2091), .Y(N33731)
         );
  NAND2BX1 U7467 ( .AN(n568), .B(n569), .Y(N34051) );
  OAI211X1 U7468 ( .A0(n7748), .A1(n1452), .B0(n2099), .C0(n2100), .Y(N33730)
         );
  OAI211X1 U7469 ( .A0(n7748), .A1(n1456), .B0(n2108), .C0(n2109), .Y(N33729)
         );
  OAI211X1 U7470 ( .A0(n7745), .A1(n1460), .B0(n2117), .C0(n2118), .Y(N33728)
         );
  NAND2BX1 U7471 ( .AN(n576), .B(n577), .Y(N34050) );
  NAND2BX1 U7472 ( .AN(n584), .B(n585), .Y(N34049) );
  NAND2BX1 U7473 ( .AN(n592), .B(n593), .Y(N34048) );
  OAI221XL U7474 ( .A0(\xArray[9][0] ), .A1(n8289), .B0(\xArray[13][0] ), .B1(
        n8235), .C0(n975), .Y(n781) );
  OAI211X1 U7475 ( .A0(n7752), .A1(n1496), .B0(n2198), .C0(n2199), .Y(N33719)
         );
  NAND2BX1 U7476 ( .AN(n664), .B(n665), .Y(N34039) );
  OAI211X1 U7477 ( .A0(n7752), .A1(n1528), .B0(n2270), .C0(n2271), .Y(N33711)
         );
  NAND2BX1 U7478 ( .AN(n728), .B(n729), .Y(N34031) );
  OAI211X1 U7479 ( .A0(n7752), .A1(n1512), .B0(n2234), .C0(n2235), .Y(N33715)
         );
  NAND2BX1 U7480 ( .AN(n696), .B(n697), .Y(N34035) );
  OAI211X1 U7481 ( .A0(n7752), .A1(n1500), .B0(n2207), .C0(n2208), .Y(N33718)
         );
  OAI211X1 U7482 ( .A0(n7752), .A1(n1504), .B0(n2216), .C0(n2217), .Y(N33717)
         );
  OAI211X1 U7483 ( .A0(n7752), .A1(n1508), .B0(n2225), .C0(n2226), .Y(N33716)
         );
  NAND2BX1 U7484 ( .AN(n672), .B(n673), .Y(N34038) );
  NAND2BX1 U7485 ( .AN(n680), .B(n681), .Y(N34037) );
  NAND2BX1 U7486 ( .AN(n688), .B(n689), .Y(N34036) );
  OAI211X1 U7487 ( .A0(n7752), .A1(n1516), .B0(n2243), .C0(n2244), .Y(N33714)
         );
  OAI211X1 U7488 ( .A0(n7752), .A1(n1520), .B0(n2252), .C0(n2253), .Y(N33713)
         );
  OAI211X1 U7489 ( .A0(n7752), .A1(n1524), .B0(n2261), .C0(n2262), .Y(N33712)
         );
  NAND2BX1 U7490 ( .AN(n704), .B(n705), .Y(N34034) );
  NAND2BX1 U7491 ( .AN(n712), .B(n713), .Y(N34033) );
  NAND2BX1 U7492 ( .AN(n720), .B(n721), .Y(N34032) );
  OAI211X1 U7493 ( .A0(n7749), .A1(n1444), .B0(n2081), .C0(n2082), .Y(N33732)
         );
  NAND2BX1 U7494 ( .AN(n560), .B(n561), .Y(N34052) );
  OAI211X1 U7495 ( .A0(n7748), .A1(n1440), .B0(n2072), .C0(n2073), .Y(N33733)
         );
  NAND2BX1 U7496 ( .AN(n552), .B(n553), .Y(N34053) );
  OAI211X1 U7497 ( .A0(n7749), .A1(n1436), .B0(n2063), .C0(n2064), .Y(N33734)
         );
  NAND2BX1 U7498 ( .AN(n544), .B(n545), .Y(N34054) );
  OAI211X1 U7499 ( .A0(n7748), .A1(n1432), .B0(n2054), .C0(n2055), .Y(N33735)
         );
  NAND2BX1 U7500 ( .AN(n536), .B(n537), .Y(N34055) );
  OAI211X1 U7501 ( .A0(n7749), .A1(n1428), .B0(n2045), .C0(n2046), .Y(N33736)
         );
  NAND2BX1 U7502 ( .AN(n528), .B(n529), .Y(N34056) );
  OAI211X1 U7503 ( .A0(n7748), .A1(n1424), .B0(n2036), .C0(n2037), .Y(N33737)
         );
  NAND2BX1 U7504 ( .AN(n520), .B(n521), .Y(N34057) );
  OAI211X1 U7505 ( .A0(n7750), .A1(n1420), .B0(n2027), .C0(n2028), .Y(N33738)
         );
  NAND2BX1 U7506 ( .AN(n512), .B(n513), .Y(N34058) );
  OAI211X1 U7507 ( .A0(n7749), .A1(n1412), .B0(n2009), .C0(n2010), .Y(N33740)
         );
  OAI211X1 U7508 ( .A0(n7744), .A1(n1416), .B0(n2018), .C0(n2019), .Y(N33739)
         );
  NAND2BX1 U7509 ( .AN(n496), .B(n497), .Y(N34060) );
  NAND2BX1 U7510 ( .AN(n504), .B(n505), .Y(N34059) );
  OAI211X1 U7511 ( .A0(n7748), .A1(n1408), .B0(n2000), .C0(n2001), .Y(N33741)
         );
  NAND2BX1 U7512 ( .AN(n488), .B(n489), .Y(N34061) );
  OAI211X1 U7513 ( .A0(n7752), .A1(n1404), .B0(n1991), .C0(n1992), .Y(N33742)
         );
  NAND2BX1 U7514 ( .AN(n480), .B(n481), .Y(N34062) );
  OAI211X1 U7515 ( .A0(n7752), .A1(n1400), .B0(n1982), .C0(n1983), .Y(N33743)
         );
  NAND2BX1 U7516 ( .AN(n472), .B(n473), .Y(N34063) );
  OAI211X1 U7517 ( .A0(n7742), .A1(n1396), .B0(n1973), .C0(n1974), .Y(N33744)
         );
  OAI211X1 U7518 ( .A0(n7742), .A1(n1392), .B0(n1964), .C0(n1965), .Y(N33745)
         );
  OAI211X1 U7519 ( .A0(n7742), .A1(n1388), .B0(n1955), .C0(n1956), .Y(N33746)
         );
  OAI211X1 U7520 ( .A0(n7742), .A1(n1384), .B0(n1946), .C0(n1947), .Y(N33747)
         );
  OAI211X1 U7521 ( .A0(n7742), .A1(n1380), .B0(n1937), .C0(n1938), .Y(N33748)
         );
  OAI211X1 U7522 ( .A0(n7742), .A1(n1376), .B0(n1928), .C0(n1929), .Y(N33749)
         );
  OAI211X1 U7523 ( .A0(n7742), .A1(n1372), .B0(n1919), .C0(n1920), .Y(N33750)
         );
  OAI211X1 U7524 ( .A0(n7742), .A1(n1368), .B0(n1910), .C0(n1911), .Y(N33751)
         );
  OAI211X1 U7525 ( .A0(n7752), .A1(n1364), .B0(n1901), .C0(n1902), .Y(N33752)
         );
  OAI211X1 U7526 ( .A0(n7744), .A1(n1360), .B0(n1892), .C0(n1893), .Y(N33753)
         );
  OAI211X1 U7527 ( .A0(n7744), .A1(n1356), .B0(n1883), .C0(n1884), .Y(N33754)
         );
  OAI211X1 U7528 ( .A0(n7746), .A1(n1352), .B0(n1874), .C0(n1875), .Y(N33755)
         );
  OAI211X1 U7529 ( .A0(n7751), .A1(n1344), .B0(n1856), .C0(n1857), .Y(N33757)
         );
  OAI211X1 U7530 ( .A0(n7751), .A1(n1348), .B0(n1865), .C0(n1866), .Y(N33756)
         );
  OAI211X1 U7531 ( .A0(n7751), .A1(n1340), .B0(n1847), .C0(n1848), .Y(N33758)
         );
  OAI211X1 U7532 ( .A0(n7751), .A1(n1336), .B0(n1838), .C0(n1839), .Y(N33759)
         );
  OAI211X1 U7533 ( .A0(n7751), .A1(n1332), .B0(n1829), .C0(n1830), .Y(N33760)
         );
  OAI211X1 U7534 ( .A0(n7751), .A1(n1328), .B0(n1820), .C0(n1821), .Y(N33761)
         );
  OAI211X1 U7535 ( .A0(n7751), .A1(n1324), .B0(n1811), .C0(n1812), .Y(N33762)
         );
  OAI211X1 U7536 ( .A0(n7751), .A1(n1320), .B0(n1802), .C0(n1803), .Y(N33763)
         );
  OAI211X1 U7537 ( .A0(n7751), .A1(n1316), .B0(n1793), .C0(n1794), .Y(N33764)
         );
  OAI211X1 U7538 ( .A0(n7751), .A1(n1312), .B0(n1784), .C0(n1785), .Y(N33765)
         );
  CLKBUFX3 U7539 ( .A(n7709), .Y(n7736) );
  OAI211X1 U7540 ( .A0(n7751), .A1(n1308), .B0(n1775), .C0(n1776), .Y(N33766)
         );
  OAI211X1 U7541 ( .A0(n7752), .A1(n1532), .B0(n2279), .C0(n2280), .Y(N33710)
         );
  OAI211X1 U7542 ( .A0(n7752), .A1(n1540), .B0(n2297), .C0(n2298), .Y(N33708)
         );
  OAI211X1 U7543 ( .A0(n7752), .A1(n1536), .B0(n2288), .C0(n2289), .Y(N33709)
         );
  NAND2BX1 U7544 ( .AN(n736), .B(n737), .Y(N34030) );
  NAND2BX1 U7545 ( .AN(n752), .B(n753), .Y(N34028) );
  NAND2BX1 U7546 ( .AN(n744), .B(n745), .Y(N34029) );
  MX4X1 U7547 ( .A(n7195), .B(n7193), .C(n7194), .D(n7192), .S0(n8407), .S1(
        N1763), .Y(N28834) );
  OAI211X1 U7548 ( .A0(n7751), .A1(n1304), .B0(n1766), .C0(n1767), .Y(N33767)
         );
  OAI221X1 U7549 ( .A0(\xArray[8][60] ), .A1(n8289), .B0(\xArray[12][60] ), 
        .B1(n8235), .C0(n993), .Y(n295) );
  CLKBUFX3 U7550 ( .A(n8221), .Y(n8218) );
  INVX3 U7551 ( .A(n8182), .Y(n8221) );
  CLKINVX1 U7552 ( .A(N1764), .Y(n6708) );
  INVX3 U7553 ( .A(n6708), .Y(n8886) );
  INVX1 U7554 ( .A(n8224), .Y(n8250) );
  CLKINVX1 U7555 ( .A(n7474), .Y(n8513) );
  CLKINVX1 U7556 ( .A(n7480), .Y(n8498) );
  INVX3 U7557 ( .A(n8306), .Y(n8334) );
  AOI221XL U7558 ( .A0(n8649), .A1(n8160), .B0(n8650), .B1(n8145), .C0(n4419), 
        .Y(n4407) );
  OAI222XL U7559 ( .A0(n8081), .A1(n3053), .B0(n8017), .B1(n3405), .C0(n8067), 
        .C1(n3124), .Y(n4419) );
  CLKINVX1 U7560 ( .A(n3336), .Y(n8647) );
  CLKINVX1 U7561 ( .A(n3541), .Y(n8646) );
  OAI222XL U7562 ( .A0(n8081), .A1(n3052), .B0(n8017), .B1(n3404), .C0(n8067), 
        .C1(n3123), .Y(n4401) );
  CLKINVX1 U7563 ( .A(n2569), .Y(n8645) );
  CLKINVX1 U7564 ( .A(n2449), .Y(n8644) );
  CLKINVX1 U7565 ( .A(n3335), .Y(n8642) );
  CLKINVX1 U7566 ( .A(n3540), .Y(n8641) );
  OAI222XL U7567 ( .A0(n8081), .A1(n3051), .B0(n8017), .B1(n3403), .C0(n8067), 
        .C1(n3122), .Y(n4383) );
  CLKINVX1 U7568 ( .A(n2568), .Y(n8640) );
  CLKINVX1 U7569 ( .A(n2446), .Y(n8639) );
  CLKINVX1 U7570 ( .A(n3334), .Y(n8637) );
  CLKINVX1 U7571 ( .A(n3539), .Y(n8636) );
  OAI222XL U7572 ( .A0(n8082), .A1(n3050), .B0(n8018), .B1(n3402), .C0(n8069), 
        .C1(n3121), .Y(n4365) );
  CLKINVX1 U7573 ( .A(n2567), .Y(n8635) );
  CLKINVX1 U7574 ( .A(n2443), .Y(n8634) );
  CLKINVX1 U7575 ( .A(n3333), .Y(n8632) );
  CLKINVX1 U7576 ( .A(n3538), .Y(n8631) );
  OAI222XL U7577 ( .A0(n8082), .A1(n3049), .B0(n8018), .B1(n3401), .C0(n8069), 
        .C1(n3120), .Y(n4347) );
  CLKINVX1 U7578 ( .A(n2566), .Y(n8630) );
  CLKINVX1 U7579 ( .A(n2440), .Y(n8629) );
  CLKINVX1 U7580 ( .A(n3332), .Y(n8627) );
  CLKINVX1 U7581 ( .A(n3537), .Y(n8626) );
  OAI222XL U7582 ( .A0(n8082), .A1(n3048), .B0(n8016), .B1(n3400), .C0(n8069), 
        .C1(n3119), .Y(n4329) );
  CLKINVX1 U7583 ( .A(n2565), .Y(n8625) );
  CLKINVX1 U7584 ( .A(n2437), .Y(n8624) );
  CLKINVX1 U7585 ( .A(n3331), .Y(n8622) );
  CLKINVX1 U7586 ( .A(n3536), .Y(n8621) );
  OAI222XL U7587 ( .A0(n8082), .A1(n3047), .B0(n8016), .B1(n3399), .C0(n8069), 
        .C1(n3118), .Y(n4311) );
  CLKINVX1 U7588 ( .A(n2564), .Y(n8620) );
  CLKINVX1 U7589 ( .A(n2434), .Y(n8619) );
  CLKINVX1 U7590 ( .A(n3330), .Y(n8617) );
  CLKINVX1 U7591 ( .A(n3535), .Y(n8616) );
  OAI222XL U7592 ( .A0(n8082), .A1(n3046), .B0(n8016), .B1(n3398), .C0(n8069), 
        .C1(n3117), .Y(n4293) );
  CLKINVX1 U7593 ( .A(n2563), .Y(n8615) );
  CLKINVX1 U7594 ( .A(n2431), .Y(n8614) );
  CLKINVX1 U7595 ( .A(n3327), .Y(n8602) );
  CLKINVX1 U7596 ( .A(n3532), .Y(n8601) );
  OAI222XL U7597 ( .A0(n8082), .A1(n3043), .B0(n8016), .B1(n3395), .C0(n8069), 
        .C1(n3114), .Y(n4239) );
  CLKINVX1 U7598 ( .A(n2560), .Y(n8600) );
  CLKINVX1 U7599 ( .A(n2422), .Y(n8599) );
  CLKINVX1 U7600 ( .A(n3326), .Y(n8597) );
  CLKINVX1 U7601 ( .A(n3531), .Y(n8596) );
  OAI222XL U7602 ( .A0(n8082), .A1(n3042), .B0(n8019), .B1(n3394), .C0(n8069), 
        .C1(n3113), .Y(n4221) );
  CLKINVX1 U7603 ( .A(n2559), .Y(n8595) );
  CLKINVX1 U7604 ( .A(n2419), .Y(n8594) );
  CLKINVX1 U7605 ( .A(n3325), .Y(n8592) );
  CLKINVX1 U7606 ( .A(n3530), .Y(n8591) );
  OAI222XL U7607 ( .A0(n8082), .A1(n3041), .B0(n6602), .B1(n3393), .C0(n8069), 
        .C1(n3112), .Y(n4203) );
  CLKINVX1 U7608 ( .A(n2558), .Y(n8590) );
  CLKINVX1 U7609 ( .A(n2416), .Y(n8589) );
  CLKINVX1 U7610 ( .A(n3324), .Y(n8587) );
  CLKINVX1 U7611 ( .A(n3529), .Y(n8586) );
  OAI222XL U7612 ( .A0(n8082), .A1(n3040), .B0(n8017), .B1(n3392), .C0(n8069), 
        .C1(n3111), .Y(n4185) );
  CLKINVX1 U7613 ( .A(n2557), .Y(n8585) );
  CLKINVX1 U7614 ( .A(n2413), .Y(n8584) );
  CLKINVX1 U7615 ( .A(n3323), .Y(n8582) );
  CLKINVX1 U7616 ( .A(n3528), .Y(n8581) );
  OAI222XL U7617 ( .A0(n8082), .A1(n3039), .B0(n8016), .B1(n3391), .C0(n8069), 
        .C1(n3110), .Y(n4167) );
  CLKINVX1 U7618 ( .A(n2556), .Y(n8580) );
  CLKINVX1 U7619 ( .A(n2410), .Y(n8579) );
  CLKINVX1 U7620 ( .A(n3322), .Y(n8577) );
  CLKINVX1 U7621 ( .A(n3527), .Y(n8576) );
  OAI222XL U7622 ( .A0(n8080), .A1(n3038), .B0(n8018), .B1(n3390), .C0(n8068), 
        .C1(n3109), .Y(n4149) );
  CLKINVX1 U7623 ( .A(n2555), .Y(n8575) );
  CLKINVX1 U7624 ( .A(n2407), .Y(n8574) );
  CLKINVX1 U7625 ( .A(n3321), .Y(n8572) );
  CLKINVX1 U7626 ( .A(n3526), .Y(n8571) );
  OAI222XL U7627 ( .A0(n8083), .A1(n3037), .B0(n8018), .B1(n3389), .C0(n8067), 
        .C1(n3108), .Y(n4131) );
  CLKINVX1 U7628 ( .A(n2554), .Y(n8570) );
  CLKINVX1 U7629 ( .A(n2404), .Y(n8569) );
  CLKINVX1 U7630 ( .A(n3320), .Y(n8567) );
  CLKINVX1 U7631 ( .A(n3525), .Y(n8566) );
  OAI222XL U7632 ( .A0(n8083), .A1(n3036), .B0(n8018), .B1(n3388), .C0(n8067), 
        .C1(n3107), .Y(n4113) );
  CLKINVX1 U7633 ( .A(n2553), .Y(n8565) );
  CLKINVX1 U7634 ( .A(n2401), .Y(n8564) );
  CLKINVX1 U7635 ( .A(n3316), .Y(n8547) );
  CLKINVX1 U7636 ( .A(n3521), .Y(n8546) );
  OAI222XL U7637 ( .A0(n8081), .A1(n3032), .B0(n8018), .B1(n3384), .C0(n8067), 
        .C1(n3103), .Y(n4041) );
  CLKINVX1 U7638 ( .A(n2549), .Y(n8545) );
  CLKINVX1 U7639 ( .A(n2389), .Y(n8544) );
  CLKINVX1 U7640 ( .A(n3315), .Y(n8542) );
  CLKINVX1 U7641 ( .A(n3520), .Y(n8541) );
  OAI222XL U7642 ( .A0(n8080), .A1(n3031), .B0(n8018), .B1(n3383), .C0(n8068), 
        .C1(n3102), .Y(n4023) );
  CLKINVX1 U7643 ( .A(n2548), .Y(n8540) );
  CLKINVX1 U7644 ( .A(n2386), .Y(n8539) );
  CLKINVX1 U7645 ( .A(n3314), .Y(n8537) );
  CLKINVX1 U7646 ( .A(n3519), .Y(n8536) );
  OAI222XL U7647 ( .A0(n8080), .A1(n3030), .B0(n8018), .B1(n3382), .C0(n8067), 
        .C1(n3101), .Y(n4005) );
  CLKINVX1 U7648 ( .A(n2547), .Y(n8535) );
  CLKINVX1 U7649 ( .A(n2383), .Y(n8534) );
  CLKINVX1 U7650 ( .A(n3311), .Y(n8522) );
  CLKINVX1 U7651 ( .A(n3516), .Y(n8521) );
  CLKINVX1 U7652 ( .A(n2544), .Y(n8520) );
  CLKINVX1 U7653 ( .A(n2374), .Y(n8519) );
  CLKINVX1 U7654 ( .A(n3313), .Y(n8532) );
  CLKINVX1 U7655 ( .A(n3518), .Y(n8531) );
  OAI222XL U7656 ( .A0(n8080), .A1(n3029), .B0(n8018), .B1(n3381), .C0(n8067), 
        .C1(n3100), .Y(n3987) );
  CLKINVX1 U7657 ( .A(n2546), .Y(n8530) );
  CLKINVX1 U7658 ( .A(n2380), .Y(n8529) );
  CLKINVX1 U7659 ( .A(n3312), .Y(n8527) );
  CLKINVX1 U7660 ( .A(n3517), .Y(n8526) );
  OAI222XL U7661 ( .A0(n8080), .A1(n3028), .B0(n8018), .B1(n3380), .C0(n8068), 
        .C1(n3099), .Y(n3969) );
  CLKINVX1 U7662 ( .A(n2545), .Y(n8525) );
  CLKINVX1 U7663 ( .A(n2377), .Y(n8524) );
  CLKINVX1 U7664 ( .A(n3309), .Y(n8512) );
  CLKINVX1 U7665 ( .A(n2368), .Y(n8509) );
  CLKINVX1 U7666 ( .A(n2542), .Y(n8510) );
  CLKINVX1 U7667 ( .A(n3308), .Y(n8507) );
  CLKINVX1 U7668 ( .A(n3513), .Y(n8506) );
  CLKINVX1 U7669 ( .A(n2365), .Y(n8504) );
  CLKINVX1 U7670 ( .A(n2541), .Y(n8505) );
  AO22X1 U7671 ( .A0(N29664), .A1(n7772), .B0(N30432), .B1(n7793), .Y(n3864)
         );
  AO22X1 U7672 ( .A0(N29667), .A1(n7773), .B0(N30435), .B1(n7793), .Y(n3810)
         );
  AO22X1 U7673 ( .A0(N29669), .A1(n7773), .B0(N30437), .B1(n7793), .Y(n3774)
         );
  CLKBUFX3 U7674 ( .A(n7710), .Y(n7739) );
  OAI22XL U7675 ( .A0(\xArray[10][56] ), .A1(n7890), .B0(n7906), .B1(n7486), 
        .Y(n3304) );
  OAI22XL U7676 ( .A0(\xArray[10][57] ), .A1(n7890), .B0(n7906), .B1(n7488), 
        .Y(n3303) );
  OAI22XL U7677 ( .A0(\xArray[10][58] ), .A1(n7890), .B0(n7907), .B1(n7490), 
        .Y(n3302) );
  OAI22XL U7678 ( .A0(\xArray[10][59] ), .A1(n7890), .B0(n7907), .B1(n7492), 
        .Y(n3301) );
  OAI22XL U7679 ( .A0(\xArray[10][61] ), .A1(n7890), .B0(n7907), .B1(n7496), 
        .Y(n3299) );
  OAI22XL U7680 ( .A0(\xArray[10][62] ), .A1(n7890), .B0(n7901), .B1(n7498), 
        .Y(n3298) );
  OAI22XL U7681 ( .A0(\xArray[7][32] ), .A1(n7848), .B0(n7859), .B1(n7439), 
        .Y(n3115) );
  OAI22XL U7682 ( .A0(\xArray[12][32] ), .A1(n7911), .B0(n7920), .B1(n7439), 
        .Y(n3465) );
  OAI22XL U7683 ( .A0(\xArray[11][32] ), .A1(n7829), .B0(n7839), .B1(n7439), 
        .Y(n3396) );
  OAI22XL U7684 ( .A0(\xArray[0][32] ), .A1(n7770), .B0(n7778), .B1(n7439), 
        .Y(n2425) );
  CLKBUFX3 U7685 ( .A(n2490), .Y(n7396) );
  CLKBUFX3 U7686 ( .A(n2487), .Y(n7398) );
  CLKBUFX3 U7687 ( .A(n2469), .Y(n7410) );
  CLKBUFX3 U7688 ( .A(n2466), .Y(n7412) );
  CLKBUFX3 U7689 ( .A(n2463), .Y(n7414) );
  OAI22XL U7690 ( .A0(\xArray[6][23] ), .A1(n7810), .B0(n7820), .B1(n7421), 
        .Y(n3053) );
  OAI22XL U7691 ( .A0(\xArray[13][24] ), .A1(n7869), .B0(n7885), .B1(n7423), 
        .Y(n3541) );
  OAI22XL U7692 ( .A0(\xArray[1][24] ), .A1(n7789), .B0(n7801), .B1(n7423), 
        .Y(n2569) );
  CLKBUFX3 U7693 ( .A(n2451), .Y(n7422) );
  OAI22XL U7694 ( .A0(\xArray[6][24] ), .A1(n7810), .B0(n7820), .B1(n7423), 
        .Y(n3052) );
  CLKBUFX3 U7695 ( .A(n2457), .Y(n7418) );
  CLKBUFX3 U7696 ( .A(n2454), .Y(n7420) );
  CLKBUFX3 U7697 ( .A(n2460), .Y(n7416) );
  CLKINVX1 U7698 ( .A(\xArray[3][1] ), .Y(n9384) );
  CLKINVX1 U7699 ( .A(\xArray[3][3] ), .Y(n9368) );
  CLKINVX1 U7700 ( .A(\xArray[3][0] ), .Y(n9392) );
  OAI22XL U7701 ( .A0(\xArray[10][49] ), .A1(n7890), .B0(n7904), .B1(n7472), 
        .Y(n3311) );
  OAI22XL U7702 ( .A0(\xArray[6][51] ), .A1(n7808), .B0(n7822), .B1(n7476), 
        .Y(n3025) );
  OAI22XL U7703 ( .A0(\xArray[10][50] ), .A1(n7890), .B0(n7905), .B1(n7474), 
        .Y(n3310) );
  OAI22XL U7704 ( .A0(\xArray[10][51] ), .A1(n7891), .B0(n7905), .B1(n7476), 
        .Y(n3309) );
  OAI22XL U7705 ( .A0(\xArray[6][52] ), .A1(n7809), .B0(n7821), .B1(n7478), 
        .Y(n3024) );
  OAI22XL U7706 ( .A0(\xArray[10][52] ), .A1(n7890), .B0(n7905), .B1(n7478), 
        .Y(n3308) );
  OAI22XL U7707 ( .A0(\xArray[10][53] ), .A1(n7890), .B0(n7905), .B1(n7480), 
        .Y(n3307) );
  OAI22XL U7708 ( .A0(\xArray[10][54] ), .A1(n7890), .B0(n7906), .B1(n7482), 
        .Y(n3306) );
  OAI22XL U7709 ( .A0(\xArray[10][55] ), .A1(n7890), .B0(n7906), .B1(n7484), 
        .Y(n3305) );
  CLKBUFX3 U7710 ( .A(n2514), .Y(n7380) );
  CLKBUFX3 U7711 ( .A(n2520), .Y(n7376) );
  CLKBUFX3 U7712 ( .A(n2517), .Y(n7378) );
  CLKBUFX3 U7713 ( .A(n2505), .Y(n7386) );
  CLKBUFX3 U7714 ( .A(n2502), .Y(n7388) );
  CLKBUFX3 U7715 ( .A(n2493), .Y(n7394) );
  CLKBUFX3 U7716 ( .A(n2511), .Y(n7382) );
  OAI22XL U7717 ( .A0(\xArray[12][24] ), .A1(n7912), .B0(n7919), .B1(n7423), 
        .Y(n3473) );
  OAI22XL U7718 ( .A0(\xArray[11][24] ), .A1(n7830), .B0(n7840), .B1(n7423), 
        .Y(n3404) );
  OAI22XL U7719 ( .A0(\xArray[12][33] ), .A1(n7911), .B0(n7920), .B1(n7441), 
        .Y(n3464) );
  OAI22XL U7720 ( .A0(\xArray[11][33] ), .A1(n7829), .B0(n7839), .B1(n7441), 
        .Y(n3395) );
  OAI22XL U7721 ( .A0(\xArray[12][35] ), .A1(n7911), .B0(n7921), .B1(n7445), 
        .Y(n3462) );
  OAI22XL U7722 ( .A0(\xArray[11][35] ), .A1(n7829), .B0(n7840), .B1(n7445), 
        .Y(n3393) );
  OAI22XL U7723 ( .A0(\xArray[12][34] ), .A1(n7911), .B0(n7921), .B1(n7443), 
        .Y(n3463) );
  OAI22XL U7724 ( .A0(\xArray[11][34] ), .A1(n7829), .B0(n7840), .B1(n7443), 
        .Y(n3394) );
  OAI22XL U7725 ( .A0(\xArray[0][35] ), .A1(n7770), .B0(n7781), .B1(n7445), 
        .Y(n2416) );
  OAI22XL U7726 ( .A0(\xArray[12][36] ), .A1(n7911), .B0(n7921), .B1(n7447), 
        .Y(n3461) );
  OAI22XL U7727 ( .A0(\xArray[11][36] ), .A1(n7829), .B0(n7840), .B1(n7447), 
        .Y(n3392) );
  OAI22XL U7728 ( .A0(\xArray[12][37] ), .A1(n7911), .B0(n7921), .B1(n7449), 
        .Y(n3460) );
  OAI22XL U7729 ( .A0(\xArray[11][37] ), .A1(n7829), .B0(n7840), .B1(n7449), 
        .Y(n3391) );
  OAI22XL U7730 ( .A0(\xArray[12][38] ), .A1(n7911), .B0(n7922), .B1(n7451), 
        .Y(n3459) );
  OAI22XL U7731 ( .A0(\xArray[11][38] ), .A1(n7829), .B0(n7841), .B1(n7451), 
        .Y(n3390) );
  OAI22XL U7732 ( .A0(\xArray[12][39] ), .A1(n7911), .B0(n7922), .B1(n7453), 
        .Y(n3458) );
  OAI22XL U7733 ( .A0(\xArray[11][39] ), .A1(n7829), .B0(n7841), .B1(n7453), 
        .Y(n3389) );
  OAI22XL U7734 ( .A0(\xArray[0][38] ), .A1(n7770), .B0(n7781), .B1(n7451), 
        .Y(n2407) );
  OAI22XL U7735 ( .A0(\xArray[7][41] ), .A1(n7851), .B0(n7860), .B1(n7457), 
        .Y(n3106) );
  OAI22XL U7736 ( .A0(\xArray[11][49] ), .A1(n7828), .B0(n7841), .B1(n7472), 
        .Y(n3379) );
  OAI22XL U7737 ( .A0(\xArray[12][49] ), .A1(n7910), .B0(n7925), .B1(n7472), 
        .Y(n3448) );
  OAI22XL U7738 ( .A0(\xArray[0][49] ), .A1(n7770), .B0(n7782), .B1(n7472), 
        .Y(n2374) );
  OAI22XL U7739 ( .A0(\xArray[11][51] ), .A1(n7828), .B0(n7841), .B1(n7476), 
        .Y(n3377) );
  OAI22XL U7740 ( .A0(\xArray[11][50] ), .A1(n7828), .B0(n7843), .B1(n7474), 
        .Y(n3378) );
  OAI22XL U7741 ( .A0(\xArray[12][50] ), .A1(n7910), .B0(n7923), .B1(n7474), 
        .Y(n3447) );
  OAI22XL U7742 ( .A0(\xArray[12][51] ), .A1(n7910), .B0(n7923), .B1(n7476), 
        .Y(n3446) );
  OAI22XL U7743 ( .A0(\xArray[0][50] ), .A1(n7769), .B0(n7779), .B1(n7474), 
        .Y(n2371) );
  OAI22XL U7744 ( .A0(\xArray[0][51] ), .A1(n7772), .B0(n7779), .B1(n7476), 
        .Y(n2368) );
  OAI22XL U7745 ( .A0(\xArray[7][51] ), .A1(n7849), .B0(n7863), .B1(n7476), 
        .Y(n3096) );
  OAI22XL U7746 ( .A0(\xArray[7][52] ), .A1(n7851), .B0(n7864), .B1(n7478), 
        .Y(n3095) );
  OAI22XL U7747 ( .A0(\xArray[11][52] ), .A1(n7828), .B0(n7843), .B1(n7478), 
        .Y(n3376) );
  OAI22XL U7748 ( .A0(\xArray[11][53] ), .A1(n7828), .B0(n7843), .B1(n7480), 
        .Y(n3375) );
  OAI22XL U7749 ( .A0(\xArray[12][52] ), .A1(n7909), .B0(n7923), .B1(n7478), 
        .Y(n3445) );
  OAI22XL U7750 ( .A0(\xArray[12][53] ), .A1(n7909), .B0(n7923), .B1(n7480), 
        .Y(n3444) );
  OAI22XL U7751 ( .A0(\xArray[0][52] ), .A1(n7773), .B0(n7778), .B1(n7478), 
        .Y(n2365) );
  OAI22XL U7752 ( .A0(\xArray[0][53] ), .A1(n7771), .B0(n7778), .B1(n7480), 
        .Y(n2362) );
  OAI22XL U7753 ( .A0(\xArray[11][54] ), .A1(n7828), .B0(n7843), .B1(n7482), 
        .Y(n3374) );
  OAI22XL U7754 ( .A0(\xArray[12][54] ), .A1(n7909), .B0(n7924), .B1(n7482), 
        .Y(n3443) );
  OAI22XL U7755 ( .A0(\xArray[0][54] ), .A1(n7771), .B0(n7781), .B1(n7482), 
        .Y(n2359) );
  OAI22XL U7756 ( .A0(\xArray[12][55] ), .A1(n7909), .B0(n7924), .B1(n7484), 
        .Y(n3442) );
  OAI22XL U7757 ( .A0(\xArray[12][56] ), .A1(n7909), .B0(n7924), .B1(n7486), 
        .Y(n3441) );
  OAI22XL U7758 ( .A0(\xArray[12][57] ), .A1(n7909), .B0(n7924), .B1(n7488), 
        .Y(n3440) );
  OAI22XL U7759 ( .A0(\xArray[12][58] ), .A1(n7909), .B0(n7925), .B1(n7490), 
        .Y(n3439) );
  OAI22XL U7760 ( .A0(\xArray[12][59] ), .A1(n7909), .B0(n7925), .B1(n7492), 
        .Y(n3438) );
  OAI22XL U7761 ( .A0(\xArray[12][61] ), .A1(n7909), .B0(n7925), .B1(n7496), 
        .Y(n3436) );
  OAI22XL U7762 ( .A0(\xArray[12][62] ), .A1(n7909), .B0(n7926), .B1(n7498), 
        .Y(n3435) );
  CLKBUFX3 U7763 ( .A(n2499), .Y(n7390) );
  CLKBUFX3 U7764 ( .A(n2496), .Y(n7392) );
  CLKBUFX3 U7765 ( .A(n2484), .Y(n7400) );
  CLKBUFX3 U7766 ( .A(n2481), .Y(n7402) );
  CLKBUFX3 U7767 ( .A(n2478), .Y(n7404) );
  CLKBUFX3 U7768 ( .A(n2472), .Y(n7408) );
  OAI22XL U7769 ( .A0(\xArray[0][24] ), .A1(n7769), .B0(n7781), .B1(n7423), 
        .Y(n2449) );
  CLKBUFX3 U7770 ( .A(n2508), .Y(n7384) );
  OAI22XL U7771 ( .A0(\xArray[0][33] ), .A1(n7770), .B0(n7774), .B1(n7441), 
        .Y(n2422) );
  OAI22XL U7772 ( .A0(\xArray[0][34] ), .A1(n7770), .B0(n7777), .B1(n7443), 
        .Y(n2419) );
  OAI22XL U7773 ( .A0(\xArray[0][36] ), .A1(n7770), .B0(n7782), .B1(n7447), 
        .Y(n2413) );
  OAI22XL U7774 ( .A0(\xArray[0][37] ), .A1(n7770), .B0(n7782), .B1(n7449), 
        .Y(n2410) );
  OAI22XL U7775 ( .A0(\xArray[12][40] ), .A1(n7910), .B0(n7922), .B1(n7455), 
        .Y(n3457) );
  OAI22XL U7776 ( .A0(\xArray[0][39] ), .A1(n7770), .B0(n7774), .B1(n7453), 
        .Y(n2404) );
  OAI22XL U7777 ( .A0(\xArray[11][40] ), .A1(n7828), .B0(n7841), .B1(n7455), 
        .Y(n3388) );
  OAI22XL U7778 ( .A0(\xArray[12][41] ), .A1(n7910), .B0(n7922), .B1(n7457), 
        .Y(n3456) );
  OAI22XL U7779 ( .A0(\xArray[11][41] ), .A1(n7828), .B0(n7841), .B1(n7457), 
        .Y(n3387) );
  OAI22XL U7780 ( .A0(\xArray[0][40] ), .A1(n7770), .B0(n7782), .B1(n7455), 
        .Y(n2401) );
  OAI22XL U7781 ( .A0(\xArray[0][41] ), .A1(n7770), .B0(n7781), .B1(n7457), 
        .Y(n2398) );
  OAI22XL U7782 ( .A0(\xArray[10][24] ), .A1(n7892), .B0(n7899), .B1(n7423), 
        .Y(n3336) );
  OAI22XL U7783 ( .A0(\xArray[6][25] ), .A1(n7810), .B0(n7820), .B1(n7425), 
        .Y(n3051) );
  OAI22XL U7784 ( .A0(\xArray[6][26] ), .A1(n7810), .B0(n7820), .B1(n7427), 
        .Y(n3050) );
  OAI22XL U7785 ( .A0(\xArray[10][25] ), .A1(n7892), .B0(n7899), .B1(n7425), 
        .Y(n3335) );
  OAI22XL U7786 ( .A0(\xArray[10][26] ), .A1(n7892), .B0(n7899), .B1(n7427), 
        .Y(n3334) );
  OAI22XL U7787 ( .A0(\xArray[6][27] ), .A1(n7810), .B0(n7821), .B1(n7429), 
        .Y(n3049) );
  OAI22XL U7788 ( .A0(\xArray[10][27] ), .A1(n7892), .B0(n7907), .B1(n7429), 
        .Y(n3333) );
  OAI22XL U7789 ( .A0(\xArray[10][28] ), .A1(n7891), .B0(n7906), .B1(n7431), 
        .Y(n3332) );
  OAI22XL U7790 ( .A0(\xArray[10][29] ), .A1(n7891), .B0(n7907), .B1(n7433), 
        .Y(n3331) );
  OAI22XL U7791 ( .A0(\xArray[10][30] ), .A1(n7891), .B0(n7906), .B1(n7435), 
        .Y(n3330) );
  OAI22XL U7792 ( .A0(\xArray[6][31] ), .A1(n7809), .B0(n7819), .B1(n7437), 
        .Y(n3045) );
  OAI22XL U7793 ( .A0(\xArray[10][31] ), .A1(n7891), .B0(n7900), .B1(n7437), 
        .Y(n3329) );
  OAI22XL U7794 ( .A0(\xArray[13][25] ), .A1(n7869), .B0(n7880), .B1(n7425), 
        .Y(n3540) );
  OAI22XL U7795 ( .A0(\xArray[1][25] ), .A1(n7789), .B0(n7801), .B1(n7425), 
        .Y(n2568) );
  OAI22XL U7796 ( .A0(\xArray[7][24] ), .A1(n7849), .B0(n7858), .B1(n7423), 
        .Y(n3123) );
  OAI22XL U7797 ( .A0(\xArray[12][25] ), .A1(n7912), .B0(n7919), .B1(n7425), 
        .Y(n3472) );
  OAI22XL U7798 ( .A0(\xArray[0][25] ), .A1(n7769), .B0(n7777), .B1(n7425), 
        .Y(n2446) );
  CLKBUFX3 U7799 ( .A(n2448), .Y(n7424) );
  AOI221XL U7800 ( .A0(n8644), .A1(n8160), .B0(n8645), .B1(n8145), .C0(n4401), 
        .Y(n4389) );
  AOI221XL U7801 ( .A0(n8646), .A1(n7993), .B0(n8647), .B1(n8030), .C0(n4398), 
        .Y(n4390) );
  OAI22XL U7802 ( .A0(\xArray[13][26] ), .A1(n7869), .B0(n7880), .B1(n7427), 
        .Y(n3539) );
  OAI22XL U7803 ( .A0(\xArray[13][27] ), .A1(n7869), .B0(n7882), .B1(n7429), 
        .Y(n3538) );
  OAI22XL U7804 ( .A0(\xArray[1][26] ), .A1(n7789), .B0(n7801), .B1(n7427), 
        .Y(n2567) );
  OAI22XL U7805 ( .A0(\xArray[1][27] ), .A1(n7789), .B0(n7800), .B1(n7429), 
        .Y(n2566) );
  OAI22XL U7806 ( .A0(\xArray[7][25] ), .A1(n7849), .B0(n7858), .B1(n7425), 
        .Y(n3122) );
  OAI22XL U7807 ( .A0(\xArray[7][26] ), .A1(n7849), .B0(n7858), .B1(n7427), 
        .Y(n3121) );
  OAI22XL U7808 ( .A0(\xArray[12][26] ), .A1(n7912), .B0(n7919), .B1(n7427), 
        .Y(n3471) );
  OAI22XL U7809 ( .A0(\xArray[12][27] ), .A1(n7912), .B0(n7921), .B1(n7429), 
        .Y(n3470) );
  OAI22XL U7810 ( .A0(\xArray[11][25] ), .A1(n7830), .B0(n7840), .B1(n7425), 
        .Y(n3403) );
  OAI22XL U7811 ( .A0(\xArray[11][26] ), .A1(n7830), .B0(n7840), .B1(n7427), 
        .Y(n3402) );
  OAI22XL U7812 ( .A0(\xArray[0][26] ), .A1(n7769), .B0(n7778), .B1(n7427), 
        .Y(n2443) );
  OAI22XL U7813 ( .A0(\xArray[0][27] ), .A1(n7769), .B0(n7777), .B1(n7429), 
        .Y(n2440) );
  CLKBUFX3 U7814 ( .A(n2445), .Y(n7426) );
  AOI221XL U7815 ( .A0(n8639), .A1(n8160), .B0(n8640), .B1(n8145), .C0(n4383), 
        .Y(n4371) );
  AOI221XL U7816 ( .A0(n8641), .A1(n7993), .B0(n8642), .B1(n8030), .C0(n4380), 
        .Y(n4372) );
  CLKBUFX3 U7817 ( .A(n2442), .Y(n7428) );
  AOI221XL U7818 ( .A0(n8634), .A1(n8160), .B0(n8635), .B1(n8145), .C0(n4365), 
        .Y(n4353) );
  AOI221XL U7819 ( .A0(n8636), .A1(n7993), .B0(n8637), .B1(n8030), .C0(n4362), 
        .Y(n4354) );
  OAI22XL U7820 ( .A0(\xArray[13][28] ), .A1(n7869), .B0(n7882), .B1(n7431), 
        .Y(n3537) );
  OAI22XL U7821 ( .A0(\xArray[13][29] ), .A1(n7869), .B0(n7883), .B1(n7433), 
        .Y(n3536) );
  OAI22XL U7822 ( .A0(\xArray[1][28] ), .A1(n7788), .B0(n7800), .B1(n7431), 
        .Y(n2565) );
  OAI22XL U7823 ( .A0(\xArray[1][29] ), .A1(n7789), .B0(n7800), .B1(n7433), 
        .Y(n2564) );
  OAI22XL U7824 ( .A0(\xArray[7][27] ), .A1(n7849), .B0(n7863), .B1(n7429), 
        .Y(n3120) );
  OAI22XL U7825 ( .A0(\xArray[12][28] ), .A1(n7911), .B0(n7922), .B1(n7431), 
        .Y(n3469) );
  OAI22XL U7826 ( .A0(\xArray[12][29] ), .A1(n7911), .B0(n7921), .B1(n7433), 
        .Y(n3468) );
  OAI22XL U7827 ( .A0(\xArray[11][27] ), .A1(n7830), .B0(n7843), .B1(n7429), 
        .Y(n3401) );
  OAI22XL U7828 ( .A0(\xArray[11][28] ), .A1(n7829), .B0(n7840), .B1(n7431), 
        .Y(n3400) );
  OAI22XL U7829 ( .A0(\xArray[0][28] ), .A1(n7769), .B0(n7777), .B1(n7431), 
        .Y(n2437) );
  OAI22XL U7830 ( .A0(\xArray[0][29] ), .A1(n7769), .B0(n7777), .B1(n7433), 
        .Y(n2434) );
  CLKBUFX3 U7831 ( .A(n2439), .Y(n7430) );
  AOI221XL U7832 ( .A0(n8629), .A1(n8160), .B0(n8630), .B1(n8145), .C0(n4347), 
        .Y(n4335) );
  AOI221XL U7833 ( .A0(n8631), .A1(n7993), .B0(n8632), .B1(n8030), .C0(n4344), 
        .Y(n4336) );
  AOI221XL U7834 ( .A0(n8624), .A1(n8160), .B0(n8625), .B1(n8145), .C0(n4329), 
        .Y(n4317) );
  AOI221XL U7835 ( .A0(n8626), .A1(n7994), .B0(n8627), .B1(n8030), .C0(n4326), 
        .Y(n4318) );
  OAI22XL U7836 ( .A0(\xArray[13][30] ), .A1(n7869), .B0(n7883), .B1(n7435), 
        .Y(n3535) );
  OAI22XL U7837 ( .A0(\xArray[13][31] ), .A1(n7870), .B0(n7882), .B1(n7437), 
        .Y(n3534) );
  OAI22XL U7838 ( .A0(\xArray[1][30] ), .A1(n7788), .B0(n7800), .B1(n7435), 
        .Y(n2563) );
  OAI22XL U7839 ( .A0(\xArray[1][31] ), .A1(n7789), .B0(n7798), .B1(n7437), 
        .Y(n2562) );
  OAI22XL U7840 ( .A0(\xArray[12][30] ), .A1(n7911), .B0(n7921), .B1(n7435), 
        .Y(n3467) );
  OAI22XL U7841 ( .A0(\xArray[12][31] ), .A1(n7911), .B0(n7920), .B1(n7437), 
        .Y(n3466) );
  OAI22XL U7842 ( .A0(\xArray[11][29] ), .A1(n7829), .B0(n7843), .B1(n7433), 
        .Y(n3399) );
  OAI22XL U7843 ( .A0(\xArray[11][30] ), .A1(n7829), .B0(n7841), .B1(n7435), 
        .Y(n3398) );
  OAI22XL U7844 ( .A0(\xArray[0][30] ), .A1(n7769), .B0(n7778), .B1(n7435), 
        .Y(n2431) );
  OAI22XL U7845 ( .A0(\xArray[0][31] ), .A1(n7770), .B0(n7777), .B1(n7437), 
        .Y(n2428) );
  CLKBUFX3 U7846 ( .A(n2433), .Y(n7434) );
  AOI221XL U7847 ( .A0(n8619), .A1(n8160), .B0(n8620), .B1(n8146), .C0(n4311), 
        .Y(n4299) );
  AOI221XL U7848 ( .A0(n8621), .A1(n7994), .B0(n8622), .B1(n8031), .C0(n4308), 
        .Y(n4300) );
  CLKBUFX3 U7849 ( .A(n2430), .Y(n7436) );
  AOI221XL U7850 ( .A0(n8614), .A1(n8160), .B0(n8615), .B1(n8146), .C0(n4293), 
        .Y(n4281) );
  AOI221XL U7851 ( .A0(n8616), .A1(n7994), .B0(n8617), .B1(n8031), .C0(n4290), 
        .Y(n4282) );
  OAI22XL U7852 ( .A0(\xArray[6][32] ), .A1(n7809), .B0(n7819), .B1(n7439), 
        .Y(n3044) );
  OAI22XL U7853 ( .A0(\xArray[10][32] ), .A1(n7891), .B0(n7900), .B1(n7439), 
        .Y(n3328) );
  OAI22XL U7854 ( .A0(\xArray[13][32] ), .A1(n7870), .B0(n7883), .B1(n7439), 
        .Y(n3533) );
  OAI22XL U7855 ( .A0(\xArray[7][31] ), .A1(n7848), .B0(n7859), .B1(n7437), 
        .Y(n3116) );
  OAI22XL U7856 ( .A0(\xArray[1][32] ), .A1(n7789), .B0(n7800), .B1(n7439), 
        .Y(n2561) );
  CLKBUFX3 U7857 ( .A(n2424), .Y(n7440) );
  AND4X1 U7858 ( .A(n4245), .B(n4246), .C(n4247), .D(n4248), .Y(n2424) );
  AOI221XL U7859 ( .A0(n7965), .A1(\xArray[9][32] ), .B0(\xArray[8][32] ), 
        .B1(n7961), .C0(n4249), .Y(n4248) );
  AOI221XL U7860 ( .A0(n8606), .A1(n7994), .B0(n8607), .B1(n8031), .C0(n4254), 
        .Y(n4246) );
  OAI22XL U7861 ( .A0(\xArray[11][31] ), .A1(n7829), .B0(n7839), .B1(n7437), 
        .Y(n3397) );
  CLKBUFX3 U7862 ( .A(n2427), .Y(n7438) );
  AND4X1 U7863 ( .A(n4263), .B(n4264), .C(n4265), .D(n4266), .Y(n2427) );
  AOI221XL U7864 ( .A0(n7965), .A1(\xArray[9][31] ), .B0(\xArray[8][31] ), 
        .B1(n7961), .C0(n4267), .Y(n4266) );
  AOI221XL U7865 ( .A0(n8611), .A1(n7994), .B0(n8612), .B1(n8031), .C0(n4272), 
        .Y(n4264) );
  OAI22XL U7866 ( .A0(\xArray[10][33] ), .A1(n7891), .B0(n7900), .B1(n7441), 
        .Y(n3327) );
  OAI22XL U7867 ( .A0(\xArray[10][34] ), .A1(n7891), .B0(n7901), .B1(n7443), 
        .Y(n3326) );
  OAI22XL U7868 ( .A0(\xArray[13][33] ), .A1(n7870), .B0(n7883), .B1(n7441), 
        .Y(n3532) );
  OAI22XL U7869 ( .A0(\xArray[13][34] ), .A1(n7870), .B0(n7883), .B1(n7443), 
        .Y(n3531) );
  OAI22XL U7870 ( .A0(\xArray[1][33] ), .A1(n7788), .B0(n7800), .B1(n7441), 
        .Y(n2560) );
  CLKBUFX3 U7871 ( .A(n2421), .Y(n7442) );
  AOI221XL U7872 ( .A0(n8599), .A1(n8160), .B0(n8600), .B1(n8146), .C0(n4239), 
        .Y(n4227) );
  AOI221XL U7873 ( .A0(n8601), .A1(n7994), .B0(n8602), .B1(n8031), .C0(n4236), 
        .Y(n4228) );
  OAI22XL U7874 ( .A0(\xArray[1][34] ), .A1(n7789), .B0(n7800), .B1(n7443), 
        .Y(n2559) );
  CLKBUFX3 U7875 ( .A(n2418), .Y(n7444) );
  AOI221XL U7876 ( .A0(n8594), .A1(n8160), .B0(n8595), .B1(n8146), .C0(n4221), 
        .Y(n4209) );
  AOI221XL U7877 ( .A0(n8596), .A1(n7994), .B0(n8597), .B1(n8031), .C0(n4218), 
        .Y(n4210) );
  OAI22XL U7878 ( .A0(\xArray[10][35] ), .A1(n7891), .B0(n7901), .B1(n7445), 
        .Y(n3325) );
  OAI22XL U7879 ( .A0(\xArray[10][36] ), .A1(n7891), .B0(n7901), .B1(n7447), 
        .Y(n3324) );
  OAI22XL U7880 ( .A0(\xArray[13][35] ), .A1(n7870), .B0(n7884), .B1(n7445), 
        .Y(n3530) );
  OAI22XL U7881 ( .A0(\xArray[13][36] ), .A1(n7870), .B0(n7883), .B1(n7447), 
        .Y(n3529) );
  OAI22XL U7882 ( .A0(\xArray[13][37] ), .A1(n7870), .B0(n7882), .B1(n7449), 
        .Y(n3528) );
  OAI22XL U7883 ( .A0(\xArray[1][35] ), .A1(n7787), .B0(n7799), .B1(n7445), 
        .Y(n2558) );
  CLKBUFX3 U7884 ( .A(n2415), .Y(n7446) );
  AOI221XL U7885 ( .A0(n8589), .A1(n8160), .B0(n8590), .B1(n8146), .C0(n4203), 
        .Y(n4191) );
  AOI221XL U7886 ( .A0(n8591), .A1(n7994), .B0(n8592), .B1(n8031), .C0(n4200), 
        .Y(n4192) );
  OAI22XL U7887 ( .A0(\xArray[1][36] ), .A1(n7788), .B0(n7799), .B1(n7447), 
        .Y(n2557) );
  CLKBUFX3 U7888 ( .A(n2412), .Y(n7448) );
  AOI221XL U7889 ( .A0(n8584), .A1(n8160), .B0(n8585), .B1(n8146), .C0(n4185), 
        .Y(n4173) );
  AOI221XL U7890 ( .A0(n8586), .A1(n7994), .B0(n8587), .B1(n8031), .C0(n4182), 
        .Y(n4174) );
  OAI22XL U7891 ( .A0(\xArray[1][37] ), .A1(n7788), .B0(n7799), .B1(n7449), 
        .Y(n2556) );
  OAI22XL U7892 ( .A0(\xArray[10][37] ), .A1(n7891), .B0(n7901), .B1(n7449), 
        .Y(n3323) );
  CLKBUFX3 U7893 ( .A(n2409), .Y(n7450) );
  AOI221XL U7894 ( .A0(n8579), .A1(n8159), .B0(n8580), .B1(n8146), .C0(n4167), 
        .Y(n4155) );
  AOI221XL U7895 ( .A0(n8581), .A1(n7994), .B0(n8582), .B1(n8031), .C0(n4164), 
        .Y(n4156) );
  OAI22XL U7896 ( .A0(\xArray[10][38] ), .A1(n7891), .B0(n7902), .B1(n7451), 
        .Y(n3322) );
  OAI22XL U7897 ( .A0(\xArray[13][38] ), .A1(n7870), .B0(n7883), .B1(n7451), 
        .Y(n3527) );
  OAI22XL U7898 ( .A0(\xArray[13][39] ), .A1(n7870), .B0(n7882), .B1(n7453), 
        .Y(n3526) );
  OAI22XL U7899 ( .A0(\xArray[1][38] ), .A1(n7787), .B0(n7799), .B1(n7451), 
        .Y(n2555) );
  CLKBUFX3 U7900 ( .A(n2406), .Y(n7452) );
  AOI221XL U7901 ( .A0(n8574), .A1(n8159), .B0(n8575), .B1(n8146), .C0(n4149), 
        .Y(n4137) );
  AOI221XL U7902 ( .A0(n8576), .A1(n7994), .B0(n8577), .B1(n8031), .C0(n4146), 
        .Y(n4138) );
  OAI22XL U7903 ( .A0(\xArray[1][39] ), .A1(n7787), .B0(n7801), .B1(n7453), 
        .Y(n2554) );
  OAI22XL U7904 ( .A0(\xArray[10][39] ), .A1(n7891), .B0(n7902), .B1(n7453), 
        .Y(n3321) );
  CLKBUFX3 U7905 ( .A(n2403), .Y(n7454) );
  AOI221XL U7906 ( .A0(n8569), .A1(n8159), .B0(n8570), .B1(n8146), .C0(n4131), 
        .Y(n4119) );
  AOI221XL U7907 ( .A0(n8571), .A1(n7994), .B0(n8572), .B1(n8031), .C0(n4128), 
        .Y(n4120) );
  OAI22XL U7908 ( .A0(\xArray[10][40] ), .A1(n7890), .B0(n7902), .B1(n7455), 
        .Y(n3320) );
  OAI22XL U7909 ( .A0(\xArray[13][40] ), .A1(n7870), .B0(n7883), .B1(n7455), 
        .Y(n3525) );
  OAI22XL U7910 ( .A0(\xArray[13][41] ), .A1(n7870), .B0(n7883), .B1(n7457), 
        .Y(n3524) );
  OAI22XL U7911 ( .A0(\xArray[1][40] ), .A1(n7788), .B0(n7798), .B1(n7455), 
        .Y(n2553) );
  CLKBUFX3 U7912 ( .A(n2400), .Y(n7456) );
  AOI221XL U7913 ( .A0(n8564), .A1(n8159), .B0(n8565), .B1(n8146), .C0(n4113), 
        .Y(n4101) );
  AOI221XL U7914 ( .A0(n8566), .A1(n7994), .B0(n8567), .B1(n8031), .C0(n4110), 
        .Y(n4102) );
  OAI22XL U7915 ( .A0(\xArray[1][41] ), .A1(n7788), .B0(n7798), .B1(n7457), 
        .Y(n2552) );
  OAI22XL U7916 ( .A0(\xArray[6][41] ), .A1(n7808), .B0(n7822), .B1(n7457), 
        .Y(n3035) );
  OAI22XL U7917 ( .A0(\xArray[6][42] ), .A1(n7808), .B0(n7821), .B1(n7459), 
        .Y(n3034) );
  OAI22XL U7918 ( .A0(\xArray[10][41] ), .A1(n7891), .B0(n7902), .B1(n7457), 
        .Y(n3319) );
  CLKBUFX3 U7919 ( .A(n2397), .Y(n7458) );
  AND4X1 U7920 ( .A(n4083), .B(n4084), .C(n4085), .D(n4086), .Y(n2397) );
  AOI221XL U7921 ( .A0(n7964), .A1(\xArray[9][41] ), .B0(\xArray[8][41] ), 
        .B1(n7960), .C0(n4087), .Y(n4086) );
  AOI221XL U7922 ( .A0(n8561), .A1(n7991), .B0(n8562), .B1(n8031), .C0(n4092), 
        .Y(n4084) );
  OAI22XL U7923 ( .A0(\xArray[10][42] ), .A1(n7891), .B0(n7903), .B1(n7459), 
        .Y(n3318) );
  OAI22XL U7924 ( .A0(\xArray[13][42] ), .A1(n7870), .B0(n7882), .B1(n7459), 
        .Y(n3523) );
  OAI22XL U7925 ( .A0(\xArray[13][43] ), .A1(n7870), .B0(n7883), .B1(n7461), 
        .Y(n3522) );
  OAI22XL U7926 ( .A0(\xArray[1][42] ), .A1(n7787), .B0(n7801), .B1(n7459), 
        .Y(n2551) );
  OAI22XL U7927 ( .A0(\xArray[1][43] ), .A1(n7787), .B0(n7802), .B1(n7461), 
        .Y(n2550) );
  OAI22XL U7928 ( .A0(\xArray[7][42] ), .A1(n7848), .B0(n7861), .B1(n7459), 
        .Y(n3105) );
  OAI22XL U7929 ( .A0(\xArray[12][42] ), .A1(n7910), .B0(n7924), .B1(n7459), 
        .Y(n3455) );
  OAI22XL U7930 ( .A0(\xArray[11][42] ), .A1(n7828), .B0(n7842), .B1(n7459), 
        .Y(n3386) );
  OAI22XL U7931 ( .A0(\xArray[12][43] ), .A1(n7910), .B0(n7926), .B1(n7461), 
        .Y(n3454) );
  OAI22XL U7932 ( .A0(\xArray[0][42] ), .A1(n7770), .B0(n7781), .B1(n7459), 
        .Y(n2395) );
  OAI22XL U7933 ( .A0(\xArray[0][43] ), .A1(n7770), .B0(n7781), .B1(n7461), 
        .Y(n2392) );
  CLKBUFX3 U7934 ( .A(n2394), .Y(n7460) );
  AND4X1 U7935 ( .A(n4065), .B(n4066), .C(n4067), .D(n4068), .Y(n2394) );
  AOI221XL U7936 ( .A0(n7964), .A1(\xArray[9][42] ), .B0(\xArray[8][42] ), 
        .B1(n7960), .C0(n4069), .Y(n4068) );
  AOI221XL U7937 ( .A0(n8556), .A1(n7991), .B0(n8557), .B1(n8031), .C0(n4074), 
        .Y(n4066) );
  OAI22XL U7938 ( .A0(\xArray[6][43] ), .A1(n7808), .B0(n7820), .B1(n7461), 
        .Y(n3033) );
  OAI22XL U7939 ( .A0(\xArray[10][43] ), .A1(n7890), .B0(n7903), .B1(n7461), 
        .Y(n3317) );
  OAI22XL U7940 ( .A0(\xArray[10][44] ), .A1(n7890), .B0(n7903), .B1(n7462), 
        .Y(n3316) );
  OAI22XL U7941 ( .A0(\xArray[13][44] ), .A1(n7871), .B0(n7883), .B1(n7462), 
        .Y(n3521) );
  OAI22XL U7942 ( .A0(\xArray[1][44] ), .A1(n7787), .B0(n7802), .B1(n7462), 
        .Y(n2549) );
  OAI22XL U7943 ( .A0(\xArray[7][43] ), .A1(n7848), .B0(n7861), .B1(n7461), 
        .Y(n3104) );
  OAI22XL U7944 ( .A0(\xArray[11][43] ), .A1(n7828), .B0(n7842), .B1(n7461), 
        .Y(n3385) );
  OAI22XL U7945 ( .A0(\xArray[12][44] ), .A1(n7910), .B0(n7921), .B1(n7462), 
        .Y(n3453) );
  OAI22XL U7946 ( .A0(\xArray[11][44] ), .A1(n7828), .B0(n7842), .B1(n7462), 
        .Y(n3384) );
  OAI22XL U7947 ( .A0(\xArray[0][44] ), .A1(n7769), .B0(n7781), .B1(n7462), 
        .Y(n2389) );
  OAI22XL U7948 ( .A0(\xArray[10][45] ), .A1(n7890), .B0(n7903), .B1(n7464), 
        .Y(n3315) );
  OAI22XL U7949 ( .A0(\xArray[10][46] ), .A1(n7890), .B0(n7904), .B1(n7466), 
        .Y(n3314) );
  OAI22XL U7950 ( .A0(\xArray[13][45] ), .A1(n7870), .B0(n7883), .B1(n7464), 
        .Y(n3520) );
  OAI22XL U7951 ( .A0(\xArray[13][46] ), .A1(n7870), .B0(n7883), .B1(n7466), 
        .Y(n3519) );
  OAI22XL U7952 ( .A0(\xArray[13][47] ), .A1(n7871), .B0(n7883), .B1(n7468), 
        .Y(n3518) );
  OAI22XL U7953 ( .A0(\xArray[1][45] ), .A1(n7787), .B0(n7799), .B1(n7464), 
        .Y(n2548) );
  OAI22XL U7954 ( .A0(\xArray[1][46] ), .A1(n7787), .B0(n7798), .B1(n7466), 
        .Y(n2547) );
  OAI22XL U7955 ( .A0(\xArray[1][47] ), .A1(n7787), .B0(n7798), .B1(n7468), 
        .Y(n2546) );
  OAI22XL U7956 ( .A0(\xArray[12][45] ), .A1(n7910), .B0(n7923), .B1(n7464), 
        .Y(n3452) );
  OAI22XL U7957 ( .A0(\xArray[11][45] ), .A1(n7828), .B0(n7842), .B1(n7464), 
        .Y(n3383) );
  OAI22XL U7958 ( .A0(\xArray[12][46] ), .A1(n7910), .B0(n7926), .B1(n7466), 
        .Y(n3451) );
  OAI22XL U7959 ( .A0(\xArray[11][46] ), .A1(n7828), .B0(n7841), .B1(n7466), 
        .Y(n3382) );
  OAI22XL U7960 ( .A0(\xArray[12][47] ), .A1(n7910), .B0(n7924), .B1(n7468), 
        .Y(n3450) );
  OAI22XL U7961 ( .A0(\xArray[11][47] ), .A1(n7828), .B0(n7841), .B1(n7468), 
        .Y(n3381) );
  CLKBUFX3 U7962 ( .A(n2388), .Y(n7463) );
  AOI221XL U7963 ( .A0(n8544), .A1(n8159), .B0(n8545), .B1(n8147), .C0(n4041), 
        .Y(n4029) );
  AOI221XL U7964 ( .A0(n8546), .A1(n7991), .B0(n8547), .B1(n8032), .C0(n4038), 
        .Y(n4030) );
  OAI22XL U7965 ( .A0(\xArray[0][45] ), .A1(n7770), .B0(n7781), .B1(n7464), 
        .Y(n2386) );
  OAI22XL U7966 ( .A0(\xArray[0][46] ), .A1(n7770), .B0(n7782), .B1(n7466), 
        .Y(n2383) );
  OAI22XL U7967 ( .A0(\xArray[0][47] ), .A1(n7769), .B0(n7781), .B1(n7468), 
        .Y(n2380) );
  CLKBUFX3 U7968 ( .A(n2385), .Y(n7465) );
  AOI221XL U7969 ( .A0(n8539), .A1(n8159), .B0(n8540), .B1(n8147), .C0(n4023), 
        .Y(n4011) );
  AOI221XL U7970 ( .A0(n8541), .A1(n7991), .B0(n8542), .B1(n8032), .C0(n4020), 
        .Y(n4012) );
  CLKBUFX3 U7971 ( .A(n2382), .Y(n7467) );
  AOI221XL U7972 ( .A0(n8534), .A1(n8159), .B0(n8535), .B1(n8147), .C0(n4005), 
        .Y(n3993) );
  AOI221XL U7973 ( .A0(n8536), .A1(n6582), .B0(n8537), .B1(n8032), .C0(n4002), 
        .Y(n3994) );
  OAI22XL U7974 ( .A0(\xArray[10][47] ), .A1(n7891), .B0(n7904), .B1(n7468), 
        .Y(n3313) );
  OAI22XL U7975 ( .A0(\xArray[10][48] ), .A1(n7891), .B0(n7904), .B1(n7470), 
        .Y(n3312) );
  OAI22XL U7976 ( .A0(\xArray[13][48] ), .A1(n7871), .B0(n7883), .B1(n7470), 
        .Y(n3517) );
  OAI22XL U7977 ( .A0(\xArray[13][49] ), .A1(n7871), .B0(n7883), .B1(n7472), 
        .Y(n3516) );
  OAI22XL U7978 ( .A0(\xArray[1][48] ), .A1(n7786), .B0(n7798), .B1(n7470), 
        .Y(n2545) );
  OAI22XL U7979 ( .A0(\xArray[1][49] ), .A1(n7786), .B0(n7798), .B1(n7472), 
        .Y(n2544) );
  CLKBUFX3 U7980 ( .A(n2373), .Y(n7473) );
  AOI221XL U7981 ( .A0(n8519), .A1(n8159), .B0(n8520), .B1(n8147), .C0(n3951), 
        .Y(n3939) );
  AOI221XL U7982 ( .A0(n8521), .A1(n7991), .B0(n8522), .B1(n8032), .C0(n3948), 
        .Y(n3940) );
  OAI22XL U7983 ( .A0(\xArray[12][48] ), .A1(n7910), .B0(n7926), .B1(n7470), 
        .Y(n3449) );
  OAI22XL U7984 ( .A0(\xArray[11][48] ), .A1(n7828), .B0(n7841), .B1(n7470), 
        .Y(n3380) );
  OAI22XL U7985 ( .A0(\xArray[0][48] ), .A1(n7769), .B0(n7782), .B1(n7470), 
        .Y(n2377) );
  CLKBUFX3 U7986 ( .A(n2379), .Y(n7469) );
  AOI221XL U7987 ( .A0(n8529), .A1(n8159), .B0(n8530), .B1(n8147), .C0(n3987), 
        .Y(n3975) );
  AOI221XL U7988 ( .A0(n8531), .A1(n7991), .B0(n8532), .B1(n8032), .C0(n3984), 
        .Y(n3976) );
  CLKBUFX3 U7989 ( .A(n2376), .Y(n7471) );
  AOI221XL U7990 ( .A0(n8524), .A1(n8159), .B0(n8525), .B1(n8147), .C0(n3969), 
        .Y(n3957) );
  AOI221XL U7991 ( .A0(n8526), .A1(n6582), .B0(n8527), .B1(n8032), .C0(n3966), 
        .Y(n3958) );
  OAI22XL U7992 ( .A0(\xArray[13][50] ), .A1(n7871), .B0(n7883), .B1(n7474), 
        .Y(n3515) );
  OAI22XL U7993 ( .A0(\xArray[13][51] ), .A1(n7871), .B0(n7883), .B1(n7476), 
        .Y(n3514) );
  OAI22XL U7994 ( .A0(\xArray[1][50] ), .A1(n7786), .B0(n7798), .B1(n7474), 
        .Y(n2543) );
  CLKBUFX3 U7995 ( .A(n2370), .Y(n7475) );
  AOI221XL U7996 ( .A0(n8514), .A1(n8159), .B0(n8515), .B1(n8147), .C0(n3933), 
        .Y(n3921) );
  OAI22XL U7997 ( .A0(\xArray[1][51] ), .A1(n7786), .B0(n7798), .B1(n7476), 
        .Y(n2542) );
  CLKBUFX3 U7998 ( .A(n2367), .Y(n7477) );
  AND4X1 U7999 ( .A(n3903), .B(n3904), .C(n3905), .D(n3906), .Y(n2367) );
  AOI221XL U8000 ( .A0(n7964), .A1(\xArray[9][51] ), .B0(\xArray[8][51] ), 
        .B1(n7960), .C0(n3907), .Y(n3906) );
  AOI221XL U8001 ( .A0(n8511), .A1(n7992), .B0(n8512), .B1(n8032), .C0(n3912), 
        .Y(n3904) );
  OAI22XL U8002 ( .A0(\xArray[13][52] ), .A1(n7871), .B0(n7882), .B1(n7478), 
        .Y(n3513) );
  OAI22XL U8003 ( .A0(\xArray[13][53] ), .A1(n7871), .B0(n7882), .B1(n7480), 
        .Y(n3512) );
  OAI22XL U8004 ( .A0(\xArray[1][52] ), .A1(n7786), .B0(n7798), .B1(n7478), 
        .Y(n2541) );
  CLKBUFX3 U8005 ( .A(n2364), .Y(n7479) );
  AND4X1 U8006 ( .A(n3885), .B(n3886), .C(n3887), .D(n3888), .Y(n2364) );
  AOI221XL U8007 ( .A0(n7963), .A1(\xArray[9][52] ), .B0(\xArray[8][52] ), 
        .B1(n7959), .C0(n3889), .Y(n3888) );
  AOI221XL U8008 ( .A0(n8506), .A1(n7991), .B0(n8507), .B1(n8032), .C0(n3894), 
        .Y(n3886) );
  OAI22XL U8009 ( .A0(\xArray[1][53] ), .A1(n7786), .B0(n7799), .B1(n7480), 
        .Y(n2540) );
  CLKBUFX3 U8010 ( .A(n2361), .Y(n7481) );
  AOI221XL U8011 ( .A0(n8499), .A1(n8158), .B0(n8500), .B1(n8147), .C0(n3879), 
        .Y(n3867) );
  OAI22XL U8012 ( .A0(\xArray[13][54] ), .A1(n7871), .B0(n7882), .B1(n7482), 
        .Y(n3511) );
  OAI22XL U8013 ( .A0(\xArray[13][55] ), .A1(n7871), .B0(n7882), .B1(n7484), 
        .Y(n3510) );
  OAI22XL U8014 ( .A0(\xArray[13][56] ), .A1(n7871), .B0(n7881), .B1(n7486), 
        .Y(n3509) );
  OAI22XL U8015 ( .A0(\xArray[1][54] ), .A1(n7786), .B0(n7798), .B1(n7482), 
        .Y(n2539) );
  CLKBUFX3 U8016 ( .A(n2358), .Y(n7483) );
  AOI221XL U8017 ( .A0(n8494), .A1(n8158), .B0(n8495), .B1(n8147), .C0(n3861), 
        .Y(n3849) );
  CLKBUFX3 U8018 ( .A(n2355), .Y(n7485) );
  AOI221XL U8019 ( .A0(n8489), .A1(n8158), .B0(n8490), .B1(n8147), .C0(n3843), 
        .Y(n3831) );
  CLKBUFX3 U8020 ( .A(n2352), .Y(n7487) );
  AOI221XL U8021 ( .A0(n8484), .A1(n8158), .B0(n8485), .B1(n8147), .C0(n3825), 
        .Y(n3813) );
  OAI22XL U8022 ( .A0(\xArray[13][57] ), .A1(n7871), .B0(n7880), .B1(n7488), 
        .Y(n3508) );
  OAI22XL U8023 ( .A0(\xArray[13][58] ), .A1(n7871), .B0(n7880), .B1(n7490), 
        .Y(n3507) );
  CLKBUFX3 U8024 ( .A(n2349), .Y(n7489) );
  AOI221XL U8025 ( .A0(n8479), .A1(n8158), .B0(n8480), .B1(n8147), .C0(n3807), 
        .Y(n3795) );
  CLKBUFX3 U8026 ( .A(n2346), .Y(n7491) );
  AOI221XL U8027 ( .A0(n8474), .A1(n8158), .B0(n8475), .B1(n8144), .C0(n3789), 
        .Y(n3777) );
  OAI22XL U8028 ( .A0(\xArray[13][59] ), .A1(n7871), .B0(n7882), .B1(n7492), 
        .Y(n3506) );
  CLKBUFX3 U8029 ( .A(n2343), .Y(n7493) );
  AOI221XL U8030 ( .A0(n8469), .A1(n8158), .B0(n8470), .B1(n8144), .C0(n3771), 
        .Y(n3759) );
  AOI221X1 U8031 ( .A0(n8464), .A1(n8158), .B0(n8465), .B1(n8146), .C0(n3753), 
        .Y(n3741) );
  OAI22XL U8032 ( .A0(\xArray[13][61] ), .A1(n7871), .B0(n7878), .B1(n7496), 
        .Y(n3504) );
  CLKBUFX3 U8033 ( .A(n2337), .Y(n7497) );
  AOI221XL U8034 ( .A0(n8454), .A1(n8158), .B0(n8455), .B1(n8144), .C0(n3735), 
        .Y(n3723) );
  OAI22XL U8035 ( .A0(\xArray[13][62] ), .A1(n7872), .B0(n7877), .B1(n7498), 
        .Y(n3503) );
  CLKBUFX3 U8036 ( .A(n2334), .Y(n7499) );
  AOI221XL U8037 ( .A0(n8449), .A1(n8158), .B0(n8450), .B1(n8145), .C0(n3717), 
        .Y(n3705) );
  CLKBUFX3 U8038 ( .A(n2328), .Y(n7501) );
  AOI221XL U8039 ( .A0(n8459), .A1(n8158), .B0(n8144), .B1(n8460), .C0(n3685), 
        .Y(n3655) );
  AOI221XL U8040 ( .A0(n6582), .A1(n8461), .B0(n8030), .B1(n8462), .C0(n3674), 
        .Y(n3656) );
  OAI221X1 U8041 ( .A0(\xArray[2][0] ), .A1(n8283), .B0(\xArray[6][0] ), .B1(
        n8229), .C0(n2323), .Y(n1742) );
  BUFX12 U8042 ( .A(n6714), .Y(n6573) );
  INVX3 U8043 ( .A(n8278), .Y(n8304) );
  CLKBUFX3 U8044 ( .A(n7707), .Y(n7732) );
  CLKBUFX3 U8045 ( .A(n7732), .Y(n7727) );
  CLKINVX3 U8046 ( .A(n8307), .Y(n8335) );
  CLKBUFX3 U8047 ( .A(n8216), .Y(n8210) );
  CLKINVX1 U8048 ( .A(n8183), .Y(n8223) );
  CLKBUFX3 U8049 ( .A(n7711), .Y(n7740) );
  INVX6 U8050 ( .A(n8327), .Y(n8314) );
  NAND2XL U8051 ( .A(n4849), .B(n773), .Y(n3689) );
  CLKBUFX2 U8052 ( .A(n8303), .Y(n8302) );
  CLKBUFX3 U8053 ( .A(n7210), .Y(n7200) );
  CLKBUFX3 U8054 ( .A(n7204), .Y(n7205) );
  CLKBUFX3 U8055 ( .A(n8410), .Y(n7210) );
  CLKBUFX3 U8056 ( .A(n7222), .Y(n7212) );
  CLKBUFX3 U8057 ( .A(n8409), .Y(n7222) );
  CLKBUFX3 U8058 ( .A(n7216), .Y(n7217) );
  NAND2XL U8059 ( .A(n4854), .B(n773), .Y(n3687) );
  AND2X1 U8060 ( .A(n8885), .B(n8886), .Y(n6574) );
  CLKBUFX3 U8061 ( .A(n7215), .Y(n7219) );
  INVX4 U8062 ( .A(n8330), .Y(n8309) );
  CLKBUFX6 U8063 ( .A(n7203), .Y(n7207) );
  INVX6 U8064 ( .A(n8328), .Y(n8312) );
  INVX3 U8065 ( .A(n8247), .Y(n8229) );
  INVX6 U8066 ( .A(n8248), .Y(n8226) );
  INVX4 U8067 ( .A(n8245), .Y(n8236) );
  INVX6 U8068 ( .A(n8304), .Y(n8283) );
  INVX4 U8069 ( .A(n8301), .Y(n8280) );
  CLKINVX1 U8070 ( .A(n6735), .Y(n266) );
  CLKBUFX3 U8071 ( .A(n6735), .Y(n8352) );
  INVX6 U8072 ( .A(n8246), .Y(n8232) );
  INVX4 U8073 ( .A(n8244), .Y(n8238) );
  INVX4 U8074 ( .A(n8248), .Y(n8241) );
  INVX6 U8075 ( .A(n8299), .Y(n8290) );
  INVX4 U8076 ( .A(n8325), .Y(n8318) );
  INVX3 U8077 ( .A(n8328), .Y(n8311) );
  NAND2X1 U8078 ( .A(n8033), .B(n8039), .Y(n6575) );
  NAND2X1 U8079 ( .A(n6611), .B(n7502), .Y(n6576) );
  NAND2X1 U8080 ( .A(n8020), .B(n8026), .Y(n6577) );
  NAND2X1 U8081 ( .A(n6619), .B(n8090), .Y(n6578) );
  NOR2X2 U8082 ( .A(n8253), .B(n7751), .Y(n6579) );
  INVX3 U8083 ( .A(n8252), .Y(n8277) );
  INVX4 U8084 ( .A(n8331), .Y(n8308) );
  INVX6 U8085 ( .A(n8245), .Y(n8235) );
  NAND2X4 U8086 ( .A(n105), .B(n106), .Y(n786) );
  CLKINVX1 U8087 ( .A(n8218), .Y(n6707) );
  INVX6 U8088 ( .A(n8300), .Y(n8286) );
  INVX4 U8089 ( .A(n8299), .Y(n8292) );
  INVX4 U8090 ( .A(n8304), .Y(n8295) );
  CLKBUFX3 U8091 ( .A(n7213), .Y(n7214) );
  NAND2X1 U8092 ( .A(n8162), .B(n8169), .Y(n6580) );
  NAND2X1 U8093 ( .A(n6617), .B(n8001), .Y(n6581) );
  NOR4X2 U8094 ( .A(n4840), .B(n6595), .C(n6601), .D(n8849), .Y(n6582) );
  BUFX2 U8095 ( .A(n8859), .Y(n7748) );
  BUFX2 U8096 ( .A(n7748), .Y(n7747) );
  BUFX2 U8097 ( .A(n8859), .Y(n7749) );
  INVX3 U8098 ( .A(n8299), .Y(n8289) );
  INVX6 U8099 ( .A(n8248), .Y(n8227) );
  INVX4 U8100 ( .A(n8324), .Y(n8323) );
  CLKBUFX3 U8101 ( .A(n7201), .Y(n7202) );
  NAND2X1 U8102 ( .A(n3293), .B(n7502), .Y(n6583) );
  NAND2X1 U8103 ( .A(n3639), .B(n7502), .Y(n6584) );
  NAND2X1 U8104 ( .A(n7992), .B(n7502), .Y(n6585) );
  NAND2X1 U8105 ( .A(n8144), .B(n7502), .Y(n6586) );
  NAND2X1 U8106 ( .A(n6615), .B(n8154), .Y(n6587) );
  NAND2X1 U8107 ( .A(n8158), .B(n7502), .Y(n6588) );
  NAND2X1 U8108 ( .A(n6618), .B(n3431), .Y(n6589) );
  NAND2X1 U8109 ( .A(n8071), .B(n3081), .Y(n6590) );
  NAND2X1 U8110 ( .A(n220), .B(n8854), .Y(n6591) );
  NAND2X1 U8111 ( .A(n181), .B(n8854), .Y(n6592) );
  NAND2X1 U8112 ( .A(n185), .B(n8854), .Y(n6593) );
  NAND2X1 U8113 ( .A(n209), .B(n8854), .Y(n6594) );
  NAND2X2 U8114 ( .A(n4831), .B(N34878), .Y(n6595) );
  NAND2X1 U8115 ( .A(n4823), .B(n8854), .Y(n6596) );
  NAND2X4 U8116 ( .A(n773), .B(n8302), .Y(n6597) );
  CLKBUFX3 U8117 ( .A(n8277), .Y(n8276) );
  NAND2X1 U8118 ( .A(n8352), .B(n8276), .Y(n1749) );
  BUFX2 U8119 ( .A(n6579), .Y(n8362) );
  BUFX4 U8120 ( .A(n7748), .Y(n7745) );
  INVX3 U8121 ( .A(n8329), .Y(n8319) );
  INVX6 U8122 ( .A(n8302), .Y(n8279) );
  INVX6 U8123 ( .A(n8249), .Y(n8225) );
  NAND2X1 U8124 ( .A(n201), .B(n8854), .Y(n6598) );
  NAND2X1 U8125 ( .A(n197), .B(n8854), .Y(n6599) );
  NAND2X1 U8126 ( .A(n205), .B(n8854), .Y(n6600) );
  NAND2X2 U8127 ( .A(n4831), .B(N34880), .Y(n6601) );
  NAND2X1 U8128 ( .A(n4859), .B(n4843), .Y(n6602) );
  OAI22X1 U8129 ( .A0(n4853), .A1(n3008), .B0(n4848), .B1(n2936), .Y(n6603) );
  AOI22X1 U8130 ( .A0(n3293), .A1(n8858), .B0(n3221), .B1(n8855), .Y(n6604) );
  CLKBUFX6 U8131 ( .A(n8178), .Y(n8177) );
  CLKBUFX6 U8132 ( .A(n8361), .Y(n8360) );
  INVX4 U8133 ( .A(n8329), .Y(n8310) );
  INVX4 U8134 ( .A(n8302), .Y(n8296) );
  INVX4 U8135 ( .A(n8249), .Y(n8242) );
  NAND2X1 U8136 ( .A(n8848), .B(n7502), .Y(n6605) );
  NAND2X1 U8137 ( .A(n8846), .B(n7502), .Y(n6606) );
  NAND2X1 U8138 ( .A(n3221), .B(n7502), .Y(n6607) );
  NAND2X1 U8139 ( .A(n2731), .B(n7502), .Y(n6608) );
  NAND2X1 U8140 ( .A(n8847), .B(n7502), .Y(n6609) );
  NOR4X2 U8141 ( .A(n4843), .B(n8850), .C(n8851), .D(n8852), .Y(n6610) );
  NOR4X2 U8142 ( .A(n6595), .B(n6601), .C(n4843), .D(n8852), .Y(n6611) );
  AND2X2 U8143 ( .A(n220), .B(n8404), .Y(n6720) );
  AND2X2 U8144 ( .A(n228), .B(n8404), .Y(n6722) );
  AND2X2 U8145 ( .A(n193), .B(n8404), .Y(n6727) );
  AND2X2 U8146 ( .A(n201), .B(n8404), .Y(n6729) );
  NAND2X1 U8147 ( .A(n232), .B(n8854), .Y(n6612) );
  NAND2X1 U8148 ( .A(n236), .B(n8854), .Y(n6613) );
  AND2X2 U8149 ( .A(n224), .B(n8404), .Y(n6721) );
  AND2X2 U8150 ( .A(n232), .B(n8404), .Y(n6723) );
  AND2X2 U8151 ( .A(n236), .B(n8404), .Y(n6724) );
  AND2X2 U8152 ( .A(n185), .B(n8404), .Y(n6725) );
  AND2X2 U8153 ( .A(n197), .B(n8404), .Y(n6728) );
  AND2X2 U8154 ( .A(n205), .B(n8404), .Y(n6730) );
  AND2X2 U8155 ( .A(n209), .B(n8404), .Y(n6731) );
  AND2X2 U8156 ( .A(n213), .B(n8404), .Y(n6732) );
  AND2X2 U8157 ( .A(n240), .B(n8404), .Y(n6733) );
  AND2X2 U8158 ( .A(n181), .B(n8404), .Y(n6734) );
  NAND2X1 U8159 ( .A(n189), .B(n8854), .Y(n6614) );
  AND2X2 U8160 ( .A(n4823), .B(n8404), .Y(n6719) );
  AND2X2 U8161 ( .A(n189), .B(n8404), .Y(n6726) );
  NOR2X1 U8162 ( .A(n8337), .B(n8279), .Y(n1747) );
  INVX6 U8163 ( .A(n8276), .Y(n8254) );
  INVX4 U8164 ( .A(n8277), .Y(n8258) );
  INVX6 U8165 ( .A(n8302), .Y(n8287) );
  INVX4 U8166 ( .A(n8201), .Y(n8198) );
  NAND2X1 U8167 ( .A(n213), .B(n8854), .Y(n6615) );
  NAND2X1 U8168 ( .A(n240), .B(n8854), .Y(n6616) );
  NAND2X1 U8169 ( .A(n224), .B(n8854), .Y(n6617) );
  NAND2X1 U8170 ( .A(n228), .B(n8854), .Y(n6618) );
  NAND2X1 U8171 ( .A(n193), .B(n8854), .Y(n6619) );
  INVX4 U8172 ( .A(n8276), .Y(n8263) );
  INVX6 U8173 ( .A(n8249), .Y(n8233) );
  CLKBUFX3 U8174 ( .A(n8179), .Y(n8181) );
  CLKBUFX2 U8175 ( .A(n3571), .Y(n7981) );
  INVX1 U8176 ( .A(n3637), .Y(n8857) );
  OAI22XL U8177 ( .A0(n7760), .A1(n782), .B0(n8350), .B1(n1292), .Y(n6621) );
  OAI22XL U8178 ( .A0(n7756), .A1(n1277), .B0(n8345), .B1(n1733), .Y(n6622) );
  AND4X4 U8179 ( .A(n4047), .B(n4048), .C(n4049), .D(n4050), .Y(n6623) );
  INVX6 U8180 ( .A(n8276), .Y(n8267) );
  CLKBUFX3 U8181 ( .A(n7750), .Y(n7741) );
  CLKBUFX3 U8182 ( .A(n8356), .Y(n8359) );
  NAND2X1 U8183 ( .A(n8352), .B(n8249), .Y(n1751) );
  CLKBUFX3 U8184 ( .A(n8170), .Y(n8172) );
  NOR2X1 U8185 ( .A(n8337), .B(n8184), .Y(n1746) );
  NOR2X1 U8186 ( .A(n8225), .B(n7751), .Y(n6714) );
  INVX6 U8187 ( .A(n8351), .Y(n8345) );
  CLKBUFX3 U8188 ( .A(n8407), .Y(n7226) );
  CLKBUFX2 U8189 ( .A(n3225), .Y(n8046) );
  CLKBUFX2 U8190 ( .A(n2942), .Y(n8097) );
  CLKBUFX2 U8191 ( .A(n2806), .Y(n8110) );
  CLKBUFX2 U8192 ( .A(n2735), .Y(n8122) );
  CLKBUFX2 U8193 ( .A(n160), .Y(n8395) );
  CLKBUFX2 U8194 ( .A(n160), .Y(n8396) );
  OAI221X4 U8195 ( .A0(n8320), .A1(n285), .B0(n7724), .B1(n791), .C0(n986), 
        .Y(N33959) );
  OAI221X4 U8196 ( .A0(n8310), .A1(n1217), .B0(n7714), .B1(n1488), .C0(n1489), 
        .Y(N33849) );
  OAI221X4 U8197 ( .A0(n8310), .A1(n1197), .B0(n7714), .B1(n1472), .C0(n1473), 
        .Y(N33853) );
  OAI221X4 U8198 ( .A0(n8310), .A1(n1177), .B0(n7714), .B1(n1456), .C0(n1457), 
        .Y(N33857) );
  OAI221X4 U8199 ( .A0(n8310), .A1(n1157), .B0(n7714), .B1(n1440), .C0(n1441), 
        .Y(N33861) );
  OAI221X4 U8200 ( .A0(n8314), .A1(n1137), .B0(n7732), .B1(n1424), .C0(n1425), 
        .Y(N33865) );
  OAI221X4 U8201 ( .A0(n8314), .A1(n1122), .B0(n7707), .B1(n1412), .C0(n1413), 
        .Y(N33868) );
  OAI221X4 U8202 ( .A0(n8314), .A1(n1107), .B0(n7712), .B1(n1400), .C0(n1401), 
        .Y(N33871) );
  OAI221X4 U8203 ( .A0(n8306), .A1(n1092), .B0(n7707), .B1(n1388), .C0(n1389), 
        .Y(N33874) );
  OAI221X4 U8204 ( .A0(n8323), .A1(n1077), .B0(n7725), .B1(n1376), .C0(n1377), 
        .Y(N33877) );
  OAI221X4 U8205 ( .A0(n8308), .A1(n1047), .B0(n7721), .B1(n1352), .C0(n1353), 
        .Y(N33883) );
  OAI221X4 U8206 ( .A0(n8308), .A1(n1032), .B0(n7711), .B1(n1340), .C0(n1341), 
        .Y(N33886) );
  OAI221X4 U8207 ( .A0(n8318), .A1(n693), .B0(n7727), .B1(n944), .C0(n1241), 
        .Y(N33908) );
  OAI221X4 U8208 ( .A0(n8319), .A1(n669), .B0(n7726), .B1(n935), .C0(n1226), 
        .Y(N33911) );
  OAI221X4 U8209 ( .A0(n8319), .A1(n645), .B0(n7726), .B1(n926), .C0(n1211), 
        .Y(N33914) );
  OAI221X4 U8210 ( .A0(n8319), .A1(n621), .B0(n7726), .B1(n917), .C0(n1196), 
        .Y(N33917) );
  OAI221X4 U8211 ( .A0(n8319), .A1(n597), .B0(n7726), .B1(n908), .C0(n1181), 
        .Y(N33920) );
  OAI221X4 U8212 ( .A0(n8320), .A1(n565), .B0(n7725), .B1(n896), .C0(n1161), 
        .Y(N33924) );
  OAI221X4 U8213 ( .A0(n8320), .A1(n517), .B0(n7725), .B1(n878), .C0(n1131), 
        .Y(N33930) );
  OAI221X4 U8214 ( .A0(n8320), .A1(n493), .B0(n7725), .B1(n869), .C0(n1116), 
        .Y(N33933) );
  OAI221X4 U8215 ( .A0(n8321), .A1(n469), .B0(n7725), .B1(n860), .C0(n1101), 
        .Y(N33936) );
  OAI221X4 U8216 ( .A0(n8321), .A1(n437), .B0(n7731), .B1(n848), .C0(n1081), 
        .Y(N33940) );
  OAI221X4 U8217 ( .A0(n8323), .A1(n413), .B0(n7731), .B1(n839), .C0(n1066), 
        .Y(N33943) );
  OAI221X4 U8218 ( .A0(n8308), .A1(n389), .B0(n7731), .B1(n830), .C0(n1051), 
        .Y(N33946) );
  OAI221X4 U8219 ( .A0(n8306), .A1(n365), .B0(n7731), .B1(n821), .C0(n1036), 
        .Y(N33949) );
  OAI221X4 U8220 ( .A0(n8308), .A1(n1052), .B0(n7725), .B1(n1356), .C0(n1357), 
        .Y(N33882) );
  OAI221X4 U8221 ( .A0(n8320), .A1(n573), .B0(n7726), .B1(n899), .C0(n1166), 
        .Y(N33923) );
  OAI221X4 U8222 ( .A0(n8314), .A1(n1132), .B0(n7732), .B1(n1420), .C0(n1421), 
        .Y(N33866) );
  OAI221X4 U8223 ( .A0(n8314), .A1(n1117), .B0(n7707), .B1(n1408), .C0(n1409), 
        .Y(N33869) );
  OAI221X4 U8224 ( .A0(n8308), .A1(n1087), .B0(n7733), .B1(n1384), .C0(n1385), 
        .Y(N33875) );
  INVX3 U8225 ( .A(n6727), .Y(n192) );
  INVX3 U8226 ( .A(n6728), .Y(n196) );
  INVX3 U8227 ( .A(n6729), .Y(n200) );
  INVX3 U8228 ( .A(n6730), .Y(n204) );
  INVX3 U8229 ( .A(n6731), .Y(n208) );
  INVX3 U8230 ( .A(n6732), .Y(n212) );
  INVX3 U8231 ( .A(n6733), .Y(n239) );
  OAI221X4 U8232 ( .A0(n8317), .A1(n767), .B0(n7723), .B1(n765), .C0(n970), 
        .Y(N33963) );
  OAI221X4 U8233 ( .A0(n8317), .A1(n751), .B0(n7723), .B1(n749), .C0(n964), 
        .Y(N33965) );
  OAI221X4 U8234 ( .A0(n8317), .A1(n759), .B0(n7723), .B1(n757), .C0(n967), 
        .Y(N33964) );
  INVX3 U8235 ( .A(n6726), .Y(n188) );
  OAI221X4 U8236 ( .A0(n8320), .A1(n293), .B0(n7724), .B1(n794), .C0(n991), 
        .Y(N33958) );
  OAI221X4 U8237 ( .A0(n8311), .A1(n1267), .B0(n7715), .B1(n1528), .C0(n1529), 
        .Y(N33839) );
  OAI221X4 U8238 ( .A0(\xArray[4][5] ), .A1(n8284), .B0(\xArray[8][5] ), .B1(
        n8230), .C0(n2278), .Y(n1528) );
  OAI221X4 U8239 ( .A0(n8320), .A1(n541), .B0(n7725), .B1(n887), .C0(n1146), 
        .Y(N33927) );
  OAI221X4 U8240 ( .A0(n8318), .A1(n701), .B0(n7727), .B1(n947), .C0(n1246), 
        .Y(N33907) );
  OAI221X4 U8241 ( .A0(n8310), .A1(n1162), .B0(n7714), .B1(n1444), .C0(n1445), 
        .Y(N33860) );
  OAI221X4 U8242 ( .A0(n8321), .A1(n445), .B0(n7731), .B1(n851), .C0(n1086), 
        .Y(N33939) );
  OAI221X4 U8243 ( .A0(n8308), .A1(n1062), .B0(n7725), .B1(n1364), .C0(n1365), 
        .Y(N33880) );
  OAI221X4 U8244 ( .A0(n8319), .A1(n589), .B0(n7726), .B1(n905), .C0(n1176), 
        .Y(N33921) );
  INVX3 U8245 ( .A(n6725), .Y(n184) );
  OAI221X4 U8246 ( .A0(n8311), .A1(n1247), .B0(n7715), .B1(n1512), .C0(n1513), 
        .Y(N33843) );
  OAI221X4 U8247 ( .A0(n8306), .A1(n317), .B0(n7724), .B1(n803), .C0(n1006), 
        .Y(N33955) );
  OAI221X4 U8248 ( .A0(n8309), .A1(n1017), .B0(n7730), .B1(n1328), .C0(n1329), 
        .Y(N33889) );
  OAI221X4 U8249 ( .A0(n8310), .A1(n1202), .B0(n7714), .B1(n1476), .C0(n1477), 
        .Y(N33852) );
  OAI221X4 U8250 ( .A0(n8323), .A1(n405), .B0(n7731), .B1(n836), .C0(n1061), 
        .Y(N33944) );
  OAI221X4 U8251 ( .A0(n8318), .A1(n717), .B0(n7727), .B1(n953), .C0(n1256), 
        .Y(N33905) );
  OAI221X4 U8252 ( .A0(\xArray[7][7] ), .A1(n8295), .B0(\xArray[11][7] ), .B1(
        n8241), .C0(n1259), .Y(n717) );
  OAI221X4 U8253 ( .A0(n8320), .A1(n509), .B0(n7725), .B1(n875), .C0(n1126), 
        .Y(N33931) );
  OAI221X4 U8254 ( .A0(n8323), .A1(n1072), .B0(n7725), .B1(n1372), .C0(n1373), 
        .Y(N33878) );
  OAI221X4 U8255 ( .A0(n8319), .A1(n613), .B0(n7726), .B1(n914), .C0(n1191), 
        .Y(N33918) );
  OAI221X4 U8256 ( .A0(n8309), .A1(n987), .B0(n7729), .B1(n1304), .C0(n1305), 
        .Y(N33895) );
  INVX3 U8257 ( .A(n6724), .Y(n235) );
  OAI221X4 U8258 ( .A0(n8311), .A1(n1232), .B0(n7715), .B1(n1500), .C0(n1501), 
        .Y(N33846) );
  OAI221X4 U8259 ( .A0(n8312), .A1(n341), .B0(n7724), .B1(n812), .C0(n1021), 
        .Y(N33952) );
  OAI221X4 U8260 ( .A0(n8314), .A1(n1102), .B0(n7711), .B1(n1396), .C0(n1397), 
        .Y(N33872) );
  OAI221X4 U8261 ( .A0(n8321), .A1(n461), .B0(n7730), .B1(n857), .C0(n1096), 
        .Y(N33937) );
  OAI221X4 U8262 ( .A0(n8309), .A1(n1027), .B0(n7711), .B1(n1336), .C0(n1337), 
        .Y(N33887) );
  OAI221X4 U8263 ( .A0(n8320), .A1(n533), .B0(n7725), .B1(n884), .C0(n1141), 
        .Y(N33928) );
  OAI221X4 U8264 ( .A0(n8310), .A1(n1172), .B0(n7714), .B1(n1452), .C0(n1453), 
        .Y(N33858) );
  OAI221X4 U8265 ( .A0(n8319), .A1(n661), .B0(n7726), .B1(n932), .C0(n1221), 
        .Y(N33912) );
  INVX3 U8266 ( .A(n6723), .Y(n231) );
  OAI221X4 U8267 ( .A0(n8309), .A1(n1002), .B0(n7711), .B1(n1316), .C0(n1317), 
        .Y(N33892) );
  OAI221X4 U8268 ( .A0(n8311), .A1(n1242), .B0(n7715), .B1(n1508), .C0(n1509), 
        .Y(N33844) );
  OAI221X4 U8269 ( .A0(n8308), .A1(n381), .B0(n7731), .B1(n827), .C0(n1046), 
        .Y(N33947) );
  OAI221X4 U8270 ( .A0(n8320), .A1(n485), .B0(n7725), .B1(n866), .C0(n1111), 
        .Y(N33934) );
  OAI221X4 U8271 ( .A0(n8312), .A1(n333), .B0(n7724), .B1(n809), .C0(n1016), 
        .Y(N33953) );
  OAI221X4 U8272 ( .A0(n8310), .A1(n1212), .B0(n7714), .B1(n1484), .C0(n1485), 
        .Y(N33850) );
  OAI221X4 U8273 ( .A0(\xArray[4][16] ), .A1(n8285), .B0(\xArray[8][16] ), 
        .B1(n8231), .C0(n2179), .Y(n1484) );
  OAI221X4 U8274 ( .A0(n8319), .A1(n637), .B0(n7726), .B1(n923), .C0(n1206), 
        .Y(N33915) );
  OAI221X4 U8275 ( .A0(n8308), .A1(n1057), .B0(n7725), .B1(n1360), .C0(n1361), 
        .Y(N33881) );
  OAI221X4 U8276 ( .A0(n8314), .A1(n1142), .B0(n7727), .B1(n1428), .C0(n1429), 
        .Y(N33864) );
  INVX3 U8277 ( .A(n6722), .Y(n227) );
  OAI221X4 U8278 ( .A0(n8311), .A1(n1257), .B0(n7715), .B1(n1520), .C0(n1521), 
        .Y(N33841) );
  OAI221X4 U8279 ( .A0(n8308), .A1(n1042), .B0(n7711), .B1(n1348), .C0(n1349), 
        .Y(N33884) );
  OAI221X4 U8280 ( .A0(n8309), .A1(n1012), .B0(n7711), .B1(n1324), .C0(n1325), 
        .Y(N33890) );
  OAI221X4 U8281 ( .A0(n8307), .A1(n357), .B0(n7724), .B1(n818), .C0(n1031), 
        .Y(N33950) );
  OAI221X4 U8282 ( .A0(n8310), .A1(n1187), .B0(n7714), .B1(n1464), .C0(n1465), 
        .Y(N33855) );
  OAI221X4 U8283 ( .A0(n8323), .A1(n421), .B0(n7731), .B1(n842), .C0(n1071), 
        .Y(N33942) );
  OAI221X4 U8284 ( .A0(n8314), .A1(n1127), .B0(n7732), .B1(n1416), .C0(n1417), 
        .Y(N33867) );
  OAI221X4 U8285 ( .A0(n8320), .A1(n525), .B0(n7725), .B1(n881), .C0(n1136), 
        .Y(N33929) );
  OAI221X4 U8286 ( .A0(n8319), .A1(n677), .B0(n7727), .B1(n938), .C0(n1231), 
        .Y(N33910) );
  INVX3 U8287 ( .A(n6721), .Y(n223) );
  OAI221X4 U8288 ( .A0(n8311), .A1(n1227), .B0(n7715), .B1(n1496), .C0(n1497), 
        .Y(N33847) );
  OAI221X4 U8289 ( .A0(n8312), .A1(n309), .B0(n7724), .B1(n800), .C0(n1001), 
        .Y(N33956) );
  OAI221X4 U8290 ( .A0(n8309), .A1(n997), .B0(n7729), .B1(n1312), .C0(n1313), 
        .Y(N33893) );
  OAI221X4 U8291 ( .A0(n8314), .A1(n1112), .B0(n7707), .B1(n1404), .C0(n1405), 
        .Y(N33870) );
  OAI221X4 U8292 ( .A0(n8318), .A1(n709), .B0(n7727), .B1(n950), .C0(n1251), 
        .Y(N33906) );
  OAI221X4 U8293 ( .A0(\xArray[7][8] ), .A1(n8295), .B0(\xArray[11][8] ), .B1(
        n8241), .C0(n1254), .Y(n709) );
  OAI221X4 U8294 ( .A0(n8308), .A1(n1037), .B0(n7711), .B1(n1344), .C0(n1345), 
        .Y(N33885) );
  OAI221X4 U8295 ( .A0(n8308), .A1(n373), .B0(n7731), .B1(n824), .C0(n1041), 
        .Y(N33948) );
  OAI221X4 U8296 ( .A0(n8320), .A1(n501), .B0(n7725), .B1(n872), .C0(n1121), 
        .Y(N33932) );
  OAI221X4 U8297 ( .A0(n8319), .A1(n605), .B0(n7726), .B1(n911), .C0(n1186), 
        .Y(N33919) );
  OAI221X4 U8298 ( .A0(n8310), .A1(n1182), .B0(n7714), .B1(n1460), .C0(n1461), 
        .Y(N33856) );
  INVX3 U8299 ( .A(n6720), .Y(n219) );
  OAI221X4 U8300 ( .A0(n8320), .A1(n397), .B0(n7731), .B1(n833), .C0(n1056), 
        .Y(N33945) );
  OAI221X4 U8301 ( .A0(n8318), .A1(n685), .B0(n7727), .B1(n941), .C0(n1236), 
        .Y(N33909) );
  OAI221X4 U8302 ( .A0(n8321), .A1(n477), .B0(n7725), .B1(n863), .C0(n1106), 
        .Y(N33935) );
  OAI221X4 U8303 ( .A0(n8314), .A1(n1097), .B0(n7711), .B1(n1392), .C0(n1393), 
        .Y(N33873) );
  OAI221X4 U8304 ( .A0(n8311), .A1(n1252), .B0(n7715), .B1(n1516), .C0(n1517), 
        .Y(N33842) );
  OAI221X4 U8305 ( .A0(\xArray[4][8] ), .A1(n8284), .B0(\xArray[8][8] ), .B1(
        n8230), .C0(n2251), .Y(n1516) );
  OAI221X4 U8306 ( .A0(n8310), .A1(n1167), .B0(n7714), .B1(n1448), .C0(n1449), 
        .Y(N33859) );
  OAI221X4 U8307 ( .A0(n8309), .A1(n1022), .B0(n7711), .B1(n1332), .C0(n1333), 
        .Y(N33888) );
  OAI221X4 U8308 ( .A0(n8307), .A1(n349), .B0(n7724), .B1(n815), .C0(n1026), 
        .Y(N33951) );
  OAI221X4 U8309 ( .A0(n8319), .A1(n581), .B0(n7726), .B1(n902), .C0(n1171), 
        .Y(N33922) );
  INVX3 U8310 ( .A(n6734), .Y(n165) );
  OAI221X4 U8311 ( .A0(n8314), .A1(n1152), .B0(n7726), .B1(n1436), .C0(n1437), 
        .Y(N33862) );
  OAI221X4 U8312 ( .A0(n8320), .A1(n557), .B0(n7725), .B1(n893), .C0(n1156), 
        .Y(N33925) );
  OAI221X4 U8313 ( .A0(n8311), .A1(n1237), .B0(n7715), .B1(n1504), .C0(n1505), 
        .Y(N33845) );
  OAI221X4 U8314 ( .A0(n8323), .A1(n1082), .B0(n7716), .B1(n1380), .C0(n1381), 
        .Y(N33876) );
  OAI221X4 U8315 ( .A0(n8321), .A1(n453), .B0(n7731), .B1(n854), .C0(n1091), 
        .Y(N33938) );
  OAI221X4 U8316 ( .A0(n8306), .A1(n325), .B0(n7724), .B1(n806), .C0(n1011), 
        .Y(N33954) );
  OAI221X4 U8317 ( .A0(n8319), .A1(n653), .B0(n7726), .B1(n929), .C0(n1216), 
        .Y(N33913) );
  OAI221X4 U8318 ( .A0(n8310), .A1(n1207), .B0(n7714), .B1(n1480), .C0(n1481), 
        .Y(N33851) );
  OAI221X4 U8319 ( .A0(n8309), .A1(n1007), .B0(n7721), .B1(n1320), .C0(n1321), 
        .Y(N33891) );
  NAND2X2 U8320 ( .A(n4831), .B(N34877), .Y(n4843) );
  NAND2X1 U8321 ( .A(n4831), .B(N34879), .Y(n4840) );
  INVX12 U8322 ( .A(n6625), .Y(x_out[31]) );
  INVX12 U8323 ( .A(n6627), .Y(x_out[30]) );
  INVX12 U8324 ( .A(n6629), .Y(x_out[29]) );
  INVX12 U8325 ( .A(n6631), .Y(x_out[28]) );
  INVX12 U8326 ( .A(n6633), .Y(x_out[27]) );
  INVX12 U8327 ( .A(n6635), .Y(x_out[26]) );
  INVX12 U8328 ( .A(n6637), .Y(x_out[25]) );
  INVX12 U8329 ( .A(n6639), .Y(x_out[24]) );
  INVX12 U8330 ( .A(n6641), .Y(x_out[23]) );
  INVX12 U8331 ( .A(n6643), .Y(x_out[22]) );
  INVX12 U8332 ( .A(n6645), .Y(x_out[21]) );
  INVX12 U8333 ( .A(n6647), .Y(x_out[20]) );
  INVX12 U8334 ( .A(n6649), .Y(x_out[19]) );
  INVX12 U8335 ( .A(n6651), .Y(x_out[18]) );
  INVX12 U8336 ( .A(n6653), .Y(x_out[17]) );
  INVX12 U8337 ( .A(n6655), .Y(x_out[16]) );
  INVX12 U8338 ( .A(n6657), .Y(x_out[15]) );
  INVX12 U8339 ( .A(n6659), .Y(x_out[14]) );
  INVX12 U8340 ( .A(n6661), .Y(x_out[13]) );
  INVX12 U8341 ( .A(n6663), .Y(x_out[12]) );
  INVX12 U8342 ( .A(n6665), .Y(x_out[11]) );
  INVX12 U8343 ( .A(n6667), .Y(x_out[10]) );
  INVX12 U8344 ( .A(n6669), .Y(x_out[9]) );
  INVX12 U8345 ( .A(n6671), .Y(x_out[8]) );
  INVX12 U8346 ( .A(n6673), .Y(x_out[7]) );
  INVX12 U8347 ( .A(n6675), .Y(x_out[6]) );
  INVX12 U8348 ( .A(n6677), .Y(x_out[5]) );
  INVX12 U8349 ( .A(n6679), .Y(x_out[4]) );
  INVX12 U8350 ( .A(n6681), .Y(x_out[3]) );
  INVX12 U8351 ( .A(n6683), .Y(x_out[2]) );
  INVX12 U8352 ( .A(n6685), .Y(x_out[1]) );
  INVX12 U8353 ( .A(n6687), .Y(x_out[0]) );
  INVX12 U8354 ( .A(n6689), .Y(out_valid) );
  INVX3 U8355 ( .A(n6719), .Y(n216) );
  OAI221X4 U8356 ( .A0(n8314), .A1(n1147), .B0(n7727), .B1(n1432), .C0(n1433), 
        .Y(N33863) );
  OAI221X4 U8357 ( .A0(n8323), .A1(n1067), .B0(n7725), .B1(n1368), .C0(n1369), 
        .Y(N33879) );
  OAI221X4 U8358 ( .A0(n8321), .A1(n429), .B0(n7731), .B1(n845), .C0(n1076), 
        .Y(N33941) );
  OAI221X4 U8359 ( .A0(n8311), .A1(n1222), .B0(n7715), .B1(n1492), .C0(n1493), 
        .Y(N33848) );
  OAI221X4 U8360 ( .A0(n8320), .A1(n549), .B0(n7725), .B1(n890), .C0(n1151), 
        .Y(N33926) );
  OAI221X4 U8361 ( .A0(n8320), .A1(n301), .B0(n7724), .B1(n797), .C0(n996), 
        .Y(N33957) );
  OAI221X4 U8362 ( .A0(n8319), .A1(n629), .B0(n7726), .B1(n920), .C0(n1201), 
        .Y(N33916) );
  OAI221X4 U8363 ( .A0(n8310), .A1(n1192), .B0(n7714), .B1(n1468), .C0(n1469), 
        .Y(N33854) );
  OAI221X4 U8364 ( .A0(n8309), .A1(n992), .B0(n7725), .B1(n1308), .C0(n1309), 
        .Y(N33894) );
  OAI221X4 U8365 ( .A0(n8318), .A1(n725), .B0(n7727), .B1(n956), .C0(n1261), 
        .Y(N33904) );
  OAI221X4 U8366 ( .A0(\xArray[7][6] ), .A1(n8295), .B0(\xArray[11][6] ), .B1(
        n8241), .C0(n1264), .Y(n725) );
  OR2X1 U8367 ( .A(\xArray[5][6] ), .B(n8281), .Y(n6691) );
  OR2X1 U8368 ( .A(\xArray[9][6] ), .B(n8227), .Y(n6692) );
  CLKINVX6 U8369 ( .A(n8301), .Y(n8281) );
  OA22X1 U8370 ( .A0(n7755), .A1(n1262), .B0(n8345), .B1(n1724), .Y(n1723) );
  OAI221X4 U8371 ( .A0(n8311), .A1(n1262), .B0(n7715), .B1(n1524), .C0(n1525), 
        .Y(N33840) );
  INVXL U8372 ( .A(n786), .Y(n6693) );
  OR2X1 U8373 ( .A(n8311), .B(n1277), .Y(n6694) );
  OR2X1 U8374 ( .A(n7715), .B(n1536), .Y(n6695) );
  NAND3X4 U8375 ( .A(n6694), .B(n6695), .C(n1537), .Y(N33837) );
  OA22X1 U8376 ( .A0(n7754), .A1(n965), .B0(n8340), .B1(n1538), .Y(n1537) );
  OR2X1 U8377 ( .A(n8318), .B(n733), .Y(n6696) );
  OR2X1 U8378 ( .A(n7727), .B(n959), .Y(n6697) );
  OAI221X4 U8379 ( .A0(\xArray[7][5] ), .A1(n8295), .B0(\xArray[11][5] ), .B1(
        n8241), .C0(n1269), .Y(n733) );
  OAI221X4 U8380 ( .A0(\xArray[6][5] ), .A1(n8292), .B0(\xArray[10][5] ), .B1(
        n8238), .C0(n1531), .Y(n959) );
  NOR2X1 U8381 ( .A(n8314), .B(n1536), .Y(n6698) );
  NOR2X1 U8382 ( .A(n7718), .B(n1538), .Y(n6699) );
  OAI221X4 U8383 ( .A0(\xArray[4][3] ), .A1(n8283), .B0(\xArray[8][3] ), .B1(
        n8229), .C0(n2296), .Y(n1536) );
  BUFX20 U8384 ( .A(n7736), .Y(n7718) );
  OAI221X4 U8385 ( .A0(\xArray[3][3] ), .A1(n8283), .B0(\xArray[7][3] ), .B1(
        n8229), .C0(n2295), .Y(n1538) );
  INVX6 U8386 ( .A(n105), .Y(n8885) );
  OAI221X4 U8387 ( .A0(n8318), .A1(n749), .B0(n7727), .B1(n965), .C0(n1276), 
        .Y(N33901) );
  INVX3 U8388 ( .A(n106), .Y(n6700) );
  OR2X1 U8389 ( .A(n8318), .B(n741), .Y(n6701) );
  OR2X1 U8390 ( .A(n7727), .B(n962), .Y(n6702) );
  OAI221X2 U8391 ( .A0(\xArray[7][4] ), .A1(n8295), .B0(\xArray[11][4] ), .B1(
        n8241), .C0(n1274), .Y(n741) );
  OAI221X4 U8392 ( .A0(\xArray[6][4] ), .A1(n8292), .B0(\xArray[10][4] ), .B1(
        n8238), .C0(n1535), .Y(n962) );
  INVX3 U8393 ( .A(n6574), .Y(n8261) );
  CLKINVX3 U8394 ( .A(n8277), .Y(n8257) );
  INVX3 U8395 ( .A(n6574), .Y(n8260) );
  CLKBUFX2 U8396 ( .A(n8218), .Y(n8206) );
  CLKINVX3 U8397 ( .A(n8300), .Y(n8284) );
  CLKINVX3 U8398 ( .A(n8246), .Y(n8230) );
  CLKBUFX2 U8399 ( .A(n6574), .Y(n8274) );
  OA22X4 U8400 ( .A0(n7756), .A1(n1282), .B0(n8345), .B1(n1736), .Y(n1735) );
  NAND3X6 U8401 ( .A(n6705), .B(n6706), .C(n1735), .Y(N33772) );
  AOI2BB2X2 U8402 ( .B0(n9382), .B1(n8207), .A0N(\xArray[10][2] ), .A1N(n8258), 
        .Y(n2302) );
  OR2X4 U8403 ( .A(\xArray[2][2] ), .B(n8283), .Y(n6703) );
  OR2X2 U8404 ( .A(\xArray[6][2] ), .B(n8229), .Y(n6704) );
  NAND3X6 U8405 ( .A(n6703), .B(n6704), .C(n2302), .Y(n1736) );
  OAI221X4 U8406 ( .A0(n8318), .A1(n757), .B0(n7727), .B1(n968), .C0(n1281), 
        .Y(N33900) );
  INVXL U8407 ( .A(n8224), .Y(n8251) );
  INVXL U8408 ( .A(n8278), .Y(n8305) );
  OA22XL U8409 ( .A0(n7760), .A1(n767), .B0(n8350), .B1(n1287), .Y(n1286) );
  OAI221X2 U8410 ( .A0(\xArray[3][2] ), .A1(n8283), .B0(\xArray[7][2] ), .B1(
        n8229), .C0(n2304), .Y(n1542) );
  OAI221X2 U8411 ( .A0(\xArray[4][2] ), .A1(n8283), .B0(\xArray[8][2] ), .B1(
        n8229), .C0(n2305), .Y(n1540) );
  INVXL U8412 ( .A(\xArray[14][2] ), .Y(n9382) );
  OA22XL U8413 ( .A0(n8323), .A1(n1542), .B0(n7728), .B1(n1736), .Y(n2297) );
  OAI221X4 U8414 ( .A0(n8318), .A1(n765), .B0(n7727), .B1(n971), .C0(n1286), 
        .Y(N33899) );
  CLKINVX2 U8415 ( .A(n7482), .Y(n8493) );
  CLKBUFX2 U8416 ( .A(n8219), .Y(n8202) );
  CLKBUFX2 U8417 ( .A(n7749), .Y(n7743) );
  OA22XL U8418 ( .A0(n7758), .A1(n758), .B0(n8347), .B1(n968), .Y(n967) );
  OA22XL U8419 ( .A0(n7756), .A1(n1272), .B0(n8345), .B1(n1730), .Y(n1729) );
  OA22XL U8420 ( .A0(n7753), .A1(n956), .B0(n8341), .B1(n1526), .Y(n1525) );
  INVX3 U8421 ( .A(n3515), .Y(n8516) );
  INVX3 U8422 ( .A(n3310), .Y(n8517) );
  NAND2XL U8423 ( .A(n8213), .B(n773), .Y(n262) );
  OA22XL U8424 ( .A0(\xArray[14][2] ), .A1(n8273), .B0(\xArray[2][2] ), .B1(
        n8187), .Y(n1543) );
  OA22XL U8425 ( .A0(\xArray[5][2] ), .A1(n8196), .B0(\xArray[1][2] ), .B1(
        n8268), .Y(n969) );
  OA22XL U8426 ( .A0(\xArray[0][6] ), .A1(n8190), .B0(\xArray[12][6] ), .B1(
        n8263), .Y(n2269) );
  OR2X1 U8427 ( .A(n8314), .B(n1540), .Y(n6705) );
  OR2X1 U8428 ( .A(n7718), .B(n1542), .Y(n6706) );
  AO22X1 U8429 ( .A0(N29661), .A1(n7772), .B0(N30429), .B1(n7793), .Y(n3918)
         );
  AO22X1 U8430 ( .A0(N29659), .A1(n7772), .B0(N30427), .B1(n7793), .Y(n3954)
         );
  AO22X1 U8431 ( .A0(N29656), .A1(n7772), .B0(N30424), .B1(n7792), .Y(n4008)
         );
  AO22X1 U8432 ( .A0(N29653), .A1(n7771), .B0(N30421), .B1(n7792), .Y(n4062)
         );
  AO22X1 U8433 ( .A0(N29648), .A1(n7771), .B0(N30416), .B1(n7792), .Y(n4152)
         );
  AO22X1 U8434 ( .A0(N29645), .A1(n7771), .B0(N30413), .B1(n7792), .Y(n4206)
         );
  AO22X1 U8435 ( .A0(N29643), .A1(n7771), .B0(N30411), .B1(n7792), .Y(n4242)
         );
  AO22X1 U8436 ( .A0(N29638), .A1(n7772), .B0(N30406), .B1(n7791), .Y(n4332)
         );
  AO22X1 U8437 ( .A0(N29640), .A1(n7771), .B0(N30408), .B1(n7792), .Y(n4296)
         );
  AO22X1 U8438 ( .A0(N29635), .A1(n7772), .B0(N30403), .B1(n7791), .Y(n4386)
         );
  AO22X1 U8439 ( .A0(N29632), .A1(n7772), .B0(N30400), .B1(n7791), .Y(n4440)
         );
  AO22X1 U8440 ( .A0(N29625), .A1(n7772), .B0(N30393), .B1(n7790), .Y(n4566)
         );
  AO22X1 U8441 ( .A0(N29623), .A1(n7772), .B0(N30391), .B1(n7790), .Y(n4602)
         );
  CLKINVX3 U8442 ( .A(n8325), .Y(n8317) );
  CLKBUFX2 U8443 ( .A(n7708), .Y(n7734) );
  NOR2XL U8444 ( .A(n8318), .B(n780), .Y(n6709) );
  NOR2XL U8445 ( .A(n7724), .B(n974), .Y(n6710) );
  OR3X6 U8446 ( .A(n6709), .B(n6710), .C(n6621), .Y(N33898) );
  NOR2X6 U8447 ( .A(n103), .B(n104), .Y(n773) );
  OAI221X1 U8448 ( .A0(\xArray[5][4] ), .A1(n8280), .B0(\xArray[9][4] ), .B1(
        n8226), .C0(n1731), .Y(n1272) );
  OAI221X4 U8449 ( .A0(n8311), .A1(n1282), .B0(n7715), .B1(n1540), .C0(n1541), 
        .Y(N33836) );
  CLKINVX2 U8450 ( .A(n7494), .Y(n8463) );
  CLKINVX2 U8451 ( .A(n7492), .Y(n8468) );
  CLKINVX2 U8452 ( .A(n7490), .Y(n8473) );
  CLKINVX2 U8453 ( .A(n7488), .Y(n8478) );
  CLKINVX2 U8454 ( .A(n7486), .Y(n8483) );
  CLKINVX2 U8455 ( .A(n7484), .Y(n8488) );
  INVX1 U8456 ( .A(n7472), .Y(n8518) );
  INVXL U8457 ( .A(n7419), .Y(n8653) );
  INVXL U8458 ( .A(n7415), .Y(n8663) );
  INVXL U8459 ( .A(n7417), .Y(n8658) );
  INVXL U8460 ( .A(n7409), .Y(n8678) );
  INVXL U8461 ( .A(n7413), .Y(n8668) );
  INVXL U8462 ( .A(n7411), .Y(n8673) );
  INVXL U8463 ( .A(n7407), .Y(n8683) );
  INVXL U8464 ( .A(n7405), .Y(n8688) );
  INVXL U8465 ( .A(n7403), .Y(n8693) );
  INVXL U8466 ( .A(n7401), .Y(n8698) );
  INVXL U8467 ( .A(n7399), .Y(n8703) );
  INVXL U8468 ( .A(n7397), .Y(n8708) );
  INVXL U8469 ( .A(n7395), .Y(n8713) );
  INVXL U8470 ( .A(n7393), .Y(n8718) );
  CLKBUFX2 U8471 ( .A(n8218), .Y(n8205) );
  CLKBUFX2 U8472 ( .A(n6574), .Y(n8275) );
  CLKBUFX2 U8473 ( .A(n7216), .Y(n7218) );
  OA22X4 U8474 ( .A0(n7756), .A1(n1292), .B0(n8345), .B1(n1742), .Y(n1741) );
  OA22XL U8475 ( .A0(n7758), .A1(n750), .B0(n8347), .B1(n965), .Y(n964) );
  OA22XL U8476 ( .A0(n7758), .A1(n742), .B0(n8347), .B1(n962), .Y(n961) );
  OA22XL U8477 ( .A0(\xArray[1][2] ), .A1(n8187), .B0(\xArray[13][2] ), .B1(
        n8260), .Y(n1737) );
  OAI221X1 U8478 ( .A0(\xArray[6][0] ), .A1(n8292), .B0(\xArray[10][0] ), .B1(
        n8238), .C0(n1551), .Y(n974) );
  NAND2X1 U8479 ( .A(n104), .B(N1761), .Y(n6711) );
  OAI221X1 U8480 ( .A0(\xArray[7][0] ), .A1(n8295), .B0(\xArray[11][0] ), .B1(
        n8241), .C0(n1294), .Y(n780) );
  INVX1 U8481 ( .A(\xArray[3][2] ), .Y(n9376) );
  OA22X2 U8482 ( .A0(\xArray[15][6] ), .A1(n8190), .B0(\xArray[11][6] ), .B1(
        n8263), .Y(n2268) );
  INVXL U8483 ( .A(\xArray[14][4] ), .Y(n9366) );
  CLKINVX3 U8484 ( .A(n8277), .Y(n8262) );
  AO22X1 U8485 ( .A0(N29630), .A1(n7772), .B0(N30398), .B1(n7791), .Y(n4476)
         );
  AO22X1 U8486 ( .A0(N29627), .A1(n7772), .B0(N30395), .B1(n7791), .Y(n4530)
         );
  CLKINVX1 U8487 ( .A(n7387), .Y(n8733) );
  CLKINVX1 U8488 ( .A(n7389), .Y(n8728) );
  CLKINVX1 U8489 ( .A(n7391), .Y(n8723) );
  AO22X1 U8490 ( .A0(N29616), .A1(n7773), .B0(N30384), .B1(n7790), .Y(n4728)
         );
  CLKINVX1 U8491 ( .A(n7381), .Y(n8748) );
  CLKINVX1 U8492 ( .A(n7383), .Y(n8743) );
  CLKINVX1 U8493 ( .A(n7385), .Y(n8738) );
  CLKINVX1 U8494 ( .A(n7375), .Y(n8763) );
  CLKINVX1 U8495 ( .A(n7377), .Y(n8758) );
  CLKINVX1 U8496 ( .A(n7379), .Y(n8753) );
  AO22X1 U8497 ( .A0(N29610), .A1(n7773), .B0(N30378), .B1(n7791), .Y(n4872)
         );
  NOR3XL U8498 ( .A(n6601), .B(n8851), .C(n4840), .Y(n4859) );
  NAND4XL U8499 ( .A(n8852), .B(n8851), .C(n8849), .D(n6601), .Y(n3080) );
  NAND4XL U8500 ( .A(n8850), .B(n4843), .C(n6595), .D(n4840), .Y(n3149) );
  OA22X2 U8501 ( .A0(n7758), .A1(n781), .B0(n8347), .B1(n974), .Y(n973) );
  OAI222XL U8502 ( .A0(n7479), .A1(n8168), .B0(n8165), .B1(n2365), .C0(n8163), 
        .C1(n7511), .Y(N28821) );
  OAI222XL U8503 ( .A0(n7477), .A1(n8168), .B0(n8165), .B1(n2368), .C0(n8163), 
        .C1(n7512), .Y(N28820) );
  OAI222XL U8504 ( .A0(n7477), .A1(n8002), .B0(n3514), .B1(n7999), .C0(n7512), 
        .C1(n7997), .Y(N27988) );
  OAI222XL U8505 ( .A0(n7477), .A1(n8041), .B0(n3309), .B1(n8037), .C0(n7512), 
        .C1(n8035), .Y(N28180) );
  OAI222XL U8506 ( .A0(n7477), .A1(n8155), .B0(n2542), .B1(n8152), .C0(n7512), 
        .C1(n8150), .Y(N28756) );
  OAI222XL U8507 ( .A0(n7479), .A1(n8002), .B0(n3513), .B1(n7998), .C0(n7511), 
        .C1(n7997), .Y(N27989) );
  OAI222XL U8508 ( .A0(n7479), .A1(n8041), .B0(n3308), .B1(n8036), .C0(n7511), 
        .C1(n8035), .Y(N28181) );
  OAI222XL U8509 ( .A0(n7479), .A1(n8155), .B0(n2541), .B1(n8151), .C0(n7511), 
        .C1(n8150), .Y(N28757) );
  OAI222XL U8510 ( .A0(n6623), .A1(n8168), .B0(n8164), .B1(n2392), .C0(n8163), 
        .C1(n7520), .Y(N28812) );
  OAI222XL U8511 ( .A0(n6623), .A1(n8002), .B0(n3522), .B1(n7999), .C0(n7520), 
        .C1(n7997), .Y(N27980) );
  OAI222XL U8512 ( .A0(n6623), .A1(n8041), .B0(n3317), .B1(n8037), .C0(n7520), 
        .C1(n8035), .Y(N28172) );
  OAI222XL U8513 ( .A0(n6623), .A1(n8155), .B0(n2550), .B1(n8152), .C0(n7520), 
        .C1(n8150), .Y(N28748) );
  OAI222XL U8514 ( .A0(n7460), .A1(n8167), .B0(n8164), .B1(n2395), .C0(n8161), 
        .C1(n7521), .Y(N28811) );
  OAI222XL U8515 ( .A0(n7458), .A1(n8001), .B0(n3524), .B1(n7999), .C0(n7522), 
        .C1(n7996), .Y(N27978) );
  OAI222XL U8516 ( .A0(n7458), .A1(n6576), .B0(n3319), .B1(n8037), .C0(n7522), 
        .C1(n8034), .Y(N28170) );
  OAI222XL U8517 ( .A0(n7458), .A1(n8156), .B0(n2552), .B1(n8152), .C0(n7522), 
        .C1(n8149), .Y(N28746) );
  OAI222XL U8518 ( .A0(n7460), .A1(n8001), .B0(n3523), .B1(n7999), .C0(n7521), 
        .C1(n7996), .Y(N27979) );
  OAI222XL U8519 ( .A0(n7460), .A1(n6576), .B0(n3318), .B1(n8037), .C0(n7521), 
        .C1(n8035), .Y(N28171) );
  OAI222XL U8520 ( .A0(n7460), .A1(n8156), .B0(n2551), .B1(n8152), .C0(n7521), 
        .C1(n8149), .Y(N28747) );
  OAI222XL U8521 ( .A0(n7438), .A1(n8167), .B0(n8166), .B1(n2428), .C0(n8161), 
        .C1(n7532), .Y(N28800) );
  OAI222XL U8522 ( .A0(n7438), .A1(n8003), .B0(n3534), .B1(n8000), .C0(n7532), 
        .C1(n7996), .Y(N27968) );
  OAI222XL U8523 ( .A0(n7438), .A1(n8041), .B0(n3329), .B1(n8038), .C0(n7532), 
        .C1(n8035), .Y(N28160) );
  OAI222XL U8524 ( .A0(n7438), .A1(n8156), .B0(n2562), .B1(n8153), .C0(n7532), 
        .C1(n8149), .Y(N28736) );
  OAI222XL U8525 ( .A0(n7440), .A1(n8003), .B0(n3533), .B1(n8000), .C0(n7531), 
        .C1(n7996), .Y(N27969) );
  OAI222XL U8526 ( .A0(n7440), .A1(n8041), .B0(n3328), .B1(n8038), .C0(n7531), 
        .C1(n8035), .Y(N28161) );
  OAI222XL U8527 ( .A0(n7440), .A1(n8156), .B0(n2561), .B1(n8153), .C0(n7531), 
        .C1(n8149), .Y(N28737) );
  AOI221XL U8528 ( .A0(n8651), .A1(n7993), .B0(n8652), .B1(n8030), .C0(n4416), 
        .Y(n4408) );
  AOI221XL U8529 ( .A0(n8696), .A1(n7993), .B0(n8697), .B1(n8030), .C0(n4578), 
        .Y(n4570) );
  AOI221XL U8530 ( .A0(n8691), .A1(n7993), .B0(n8692), .B1(n8030), .C0(n4560), 
        .Y(n4552) );
  AOI221XL U8531 ( .A0(n8686), .A1(n7993), .B0(n8687), .B1(n8030), .C0(n4542), 
        .Y(n4534) );
  AOI221XL U8532 ( .A0(n8681), .A1(n7993), .B0(n8682), .B1(n8030), .C0(n4524), 
        .Y(n4516) );
  AOI221XL U8533 ( .A0(n8701), .A1(n7992), .B0(n8702), .B1(n6611), .C0(n4596), 
        .Y(n4588) );
  AOI221XL U8534 ( .A0(n8731), .A1(n7992), .B0(n8732), .B1(n6611), .C0(n4704), 
        .Y(n4696) );
  AOI221XL U8535 ( .A0(n8726), .A1(n7992), .B0(n8727), .B1(n8029), .C0(n4686), 
        .Y(n4678) );
  AOI221XL U8536 ( .A0(n8721), .A1(n7992), .B0(n8722), .B1(n8029), .C0(n4668), 
        .Y(n4660) );
  AOI221XL U8537 ( .A0(n8716), .A1(n7992), .B0(n8717), .B1(n8029), .C0(n4650), 
        .Y(n4642) );
  AOI221XL U8538 ( .A0(n8746), .A1(n7992), .B0(n8747), .B1(n8029), .C0(n4758), 
        .Y(n4750) );
  AOI221XL U8539 ( .A0(n8741), .A1(n7992), .B0(n8742), .B1(n8029), .C0(n4740), 
        .Y(n4732) );
  AOI221XL U8540 ( .A0(n8736), .A1(n7992), .B0(n8737), .B1(n8029), .C0(n4722), 
        .Y(n4714) );
  AOI221XL U8541 ( .A0(n8756), .A1(n7992), .B0(n8757), .B1(n8029), .C0(n4794), 
        .Y(n4786) );
  AOI221XL U8542 ( .A0(n8751), .A1(n7992), .B0(n8752), .B1(n8029), .C0(n4776), 
        .Y(n4768) );
  NAND2XL U8543 ( .A(n4883), .B(n216), .Y(N1805) );
  OAI221X1 U8544 ( .A0(\xArray[4][4] ), .A1(n8283), .B0(\xArray[8][4] ), .B1(
        n8229), .C0(n2287), .Y(n1532) );
  AOI2BB2XL U8545 ( .B0(n9390), .B1(n8207), .A0N(\xArray[10][1] ), .A1N(n8258), 
        .Y(n2311) );
  OA22XL U8546 ( .A0(\xArray[14][4] ), .A1(n8272), .B0(\xArray[2][4] ), .B1(
        n8186), .Y(n1535) );
  INVX1 U8547 ( .A(\xArray[14][5] ), .Y(n9358) );
  INVXL U8548 ( .A(\xArray[14][0] ), .Y(n9398) );
  INVX1 U8549 ( .A(\xArray[14][6] ), .Y(n9350) );
  INVXL U8550 ( .A(\xArray[14][1] ), .Y(n9390) );
  MX4X1 U8551 ( .A(\bArray[0][34] ), .B(\bArray[1][34] ), .C(\bArray[2][34] ), 
        .D(\bArray[3][34] ), .S0(n7201), .S1(N1762), .Y(n7083) );
  CLKINVX1 U8552 ( .A(\xArray[14][38] ), .Y(n9094) );
  CLKINVX1 U8553 ( .A(\xArray[14][39] ), .Y(n9086) );
  CLKINVX1 U8554 ( .A(\xArray[14][40] ), .Y(n9078) );
  INVX1 U8555 ( .A(n6711), .Y(n2325) );
  OR2X1 U8556 ( .A(n8311), .B(n1272), .Y(n6712) );
  OR2XL U8557 ( .A(n7715), .B(n1532), .Y(n6713) );
  NAND3X4 U8558 ( .A(n6712), .B(n6713), .C(n1533), .Y(N33838) );
  OA22XL U8559 ( .A0(n7753), .A1(n962), .B0(n8340), .B1(n1534), .Y(n1533) );
  CLKBUFX2 U8560 ( .A(n8362), .Y(n8361) );
  CLKBUFX2 U8561 ( .A(n8176), .Y(n8178) );
  CLKINVX3 U8562 ( .A(n8276), .Y(n8259) );
  CLKINVX3 U8563 ( .A(n8277), .Y(n8264) );
  INVX1 U8564 ( .A(n7478), .Y(n8503) );
  INVX1 U8565 ( .A(n7476), .Y(n8508) );
  CLKINVX3 U8566 ( .A(n8276), .Y(n8255) );
  INVX1 U8567 ( .A(n7470), .Y(n8523) );
  INVX1 U8568 ( .A(n7468), .Y(n8528) );
  CLKINVX3 U8569 ( .A(n8277), .Y(n8265) );
  INVX1 U8570 ( .A(n7466), .Y(n8533) );
  INVX1 U8571 ( .A(n7464), .Y(n8538) );
  INVX1 U8572 ( .A(n7462), .Y(n8543) );
  INVX1 U8573 ( .A(n7461), .Y(n8548) );
  INVX1 U8574 ( .A(n7459), .Y(n8553) );
  INVX1 U8575 ( .A(n7457), .Y(n8558) );
  INVX1 U8576 ( .A(n7455), .Y(n8563) );
  INVX1 U8577 ( .A(n7453), .Y(n8568) );
  INVX1 U8578 ( .A(n7451), .Y(n8573) );
  CLKINVX3 U8579 ( .A(n8276), .Y(n8266) );
  INVX1 U8580 ( .A(n7449), .Y(n8578) );
  INVX1 U8581 ( .A(n7447), .Y(n8583) );
  INVX1 U8582 ( .A(n7445), .Y(n8588) );
  INVX1 U8583 ( .A(n7443), .Y(n8593) );
  INVX1 U8584 ( .A(n7441), .Y(n8598) );
  INVX1 U8585 ( .A(n7435), .Y(n8613) );
  INVX1 U8586 ( .A(n7439), .Y(n8603) );
  INVX1 U8587 ( .A(n7437), .Y(n8608) );
  INVX1 U8588 ( .A(n7433), .Y(n8618) );
  INVX1 U8589 ( .A(n7431), .Y(n8623) );
  INVX1 U8590 ( .A(n7429), .Y(n8628) );
  CLKINVX3 U8591 ( .A(n8276), .Y(n8256) );
  INVX1 U8592 ( .A(n7427), .Y(n8633) );
  INVX1 U8593 ( .A(n7425), .Y(n8638) );
  INVX1 U8594 ( .A(n7423), .Y(n8643) );
  INVX1 U8595 ( .A(n7421), .Y(n8648) );
  INVX3 U8596 ( .A(n7796), .Y(n7791) );
  INVX3 U8597 ( .A(n7795), .Y(n7792) );
  BUFX12 U8598 ( .A(n2600), .Y(n7500) );
  AOI221X2 U8599 ( .A0(N33705), .A1(n7875), .B0(N31401), .B1(n7700), .C0(n3699), .Y(n3697) );
  BUFX12 U8600 ( .A(n2605), .Y(n7496) );
  AOI221X2 U8601 ( .A0(N33703), .A1(n7874), .B0(N31399), .B1(n7703), .C0(n3738), .Y(n3737) );
  BUFX12 U8602 ( .A(n2603), .Y(n7498) );
  AOI221X2 U8603 ( .A0(N33704), .A1(n7875), .B0(N31400), .B1(n7703), .C0(n3720), .Y(n3719) );
  CLKBUFX2 U8604 ( .A(n8218), .Y(n8207) );
  AO22X4 U8605 ( .A0(N29670), .A1(n7773), .B0(N30438), .B1(n7793), .Y(n3756)
         );
  CLKINVX3 U8606 ( .A(n8299), .Y(n8293) );
  CLKINVX3 U8607 ( .A(n8244), .Y(n8239) );
  CLKINVX3 U8608 ( .A(n8300), .Y(n8285) );
  CLKINVX3 U8609 ( .A(n8246), .Y(n8231) );
  CLKINVX3 U8610 ( .A(n8325), .Y(n8316) );
  CLKBUFX2 U8611 ( .A(n8217), .Y(n8209) );
  CLKINVX3 U8612 ( .A(n8327), .Y(n8313) );
  CLKINVX3 U8613 ( .A(n8302), .Y(n8297) );
  CLKINVX3 U8614 ( .A(n8249), .Y(n8243) );
  CLKINVX2 U8615 ( .A(n8324), .Y(n8322) );
  CLKBUFX2 U8616 ( .A(n8219), .Y(n8203) );
  CLKINVX3 U8617 ( .A(n8245), .Y(n8237) );
  CLKINVX3 U8618 ( .A(n8299), .Y(n8291) );
  CLKINVX3 U8619 ( .A(n8302), .Y(n8282) );
  CLKINVX3 U8620 ( .A(n8247), .Y(n8228) );
  CLKINVX3 U8621 ( .A(n8302), .Y(n8294) );
  CLKINVX3 U8622 ( .A(n8249), .Y(n8240) );
  CLKINVX3 U8623 ( .A(n8302), .Y(n8288) );
  CLKINVX3 U8624 ( .A(n8249), .Y(n8234) );
  CLKINVX3 U8625 ( .A(n8332), .Y(n8320) );
  CLKINVX2 U8626 ( .A(n8302), .Y(n8298) );
  CLKINVX2 U8627 ( .A(n8201), .Y(n8200) );
  CLKINVX3 U8628 ( .A(n8201), .Y(n8199) );
  CLKBUFX3 U8629 ( .A(n8856), .Y(n7700) );
  CLKBUFX3 U8630 ( .A(n8857), .Y(n7705) );
  CLKBUFX3 U8631 ( .A(n8857), .Y(n7706) );
  CLKBUFX3 U8632 ( .A(n8856), .Y(n7701) );
  CLKBUFX3 U8633 ( .A(n8856), .Y(n7702) );
  CLKBUFX3 U8634 ( .A(n7736), .Y(n7719) );
  BUFX8 U8635 ( .A(n7708), .Y(n7735) );
  CLKBUFX2 U8636 ( .A(n7710), .Y(n7738) );
  CLKBUFX2 U8637 ( .A(n7749), .Y(n7744) );
  CLKBUFX2 U8638 ( .A(n7748), .Y(n7746) );
  CLKBUFX2 U8639 ( .A(n7750), .Y(n7742) );
  CLKBUFX2 U8640 ( .A(n8215), .Y(n8212) );
  CLKBUFX2 U8641 ( .A(n7708), .Y(n7733) );
  CLKBUFX2 U8642 ( .A(n7709), .Y(n7737) );
  CLKINVX3 U8643 ( .A(n8351), .Y(n8344) );
  CLKINVX3 U8644 ( .A(n8351), .Y(n8346) );
  CLKINVX3 U8645 ( .A(n8352), .Y(n8349) );
  CLKBUFX2 U8646 ( .A(n7707), .Y(n7731) );
  CLKBUFX2 U8647 ( .A(n7215), .Y(n7220) );
  CLKBUFX2 U8648 ( .A(n8356), .Y(n8358) );
  CLKINVX3 U8649 ( .A(n8351), .Y(n8343) );
  CLKINVX3 U8650 ( .A(n8352), .Y(n8348) );
  CLKINVX1 U8651 ( .A(N25664), .Y(n8768) );
  AND2X2 U8652 ( .A(n2728), .B(n2729), .Y(n2601) );
  AND2X2 U8653 ( .A(n3218), .B(n3219), .Y(n3154) );
  CLKINVX1 U8654 ( .A(n2729), .Y(n8856) );
  OR2X1 U8655 ( .A(n4833), .B(n7761), .Y(n3662) );
  INVX1 U8656 ( .A(n8278), .Y(n8303) );
  INVXL U8657 ( .A(n8182), .Y(n8222) );
  INVXL U8658 ( .A(n8306), .Y(n8333) );
  INVXL U8659 ( .A(n8307), .Y(n8336) );
  NAND2XL U8660 ( .A(n4861), .B(n8352), .Y(n3695) );
  INVX1 U8661 ( .A(n6595), .Y(n8851) );
  NAND2X1 U8662 ( .A(n4858), .B(n8332), .Y(n3637) );
  CLKINVX1 U8663 ( .A(n4843), .Y(n8849) );
  CLKINVX1 U8664 ( .A(n4822), .Y(n8860) );
  NAND2XL U8665 ( .A(n4849), .B(n8352), .Y(n3219) );
  NAND2XL U8666 ( .A(n4858), .B(n8352), .Y(n3678) );
  INVX3 U8667 ( .A(n2331), .Y(n8459) );
  INVX3 U8668 ( .A(n2528), .Y(n8460) );
  OAI222X2 U8669 ( .A0(n3011), .A1(n8080), .B0(n3363), .B1(n8016), .C0(n3082), 
        .C1(n8068), .Y(n3685) );
  INVX3 U8670 ( .A(n2338), .Y(n8454) );
  INVX3 U8671 ( .A(n2532), .Y(n8455) );
  OAI222X2 U8672 ( .A0(n8083), .A1(n3015), .B0(n8019), .B1(n3367), .C0(n8070), 
        .C1(n3086), .Y(n3735) );
  INVX3 U8673 ( .A(n2335), .Y(n8449) );
  INVX3 U8674 ( .A(n2531), .Y(n8450) );
  INVX3 U8675 ( .A(n2341), .Y(n8464) );
  INVX3 U8676 ( .A(n2533), .Y(n8465) );
  OAI222X2 U8677 ( .A0(n8083), .A1(n3016), .B0(n8019), .B1(n3368), .C0(n8070), 
        .C1(n3087), .Y(n3753) );
  AOI221X2 U8678 ( .A0(n8456), .A1(n7991), .B0(n8457), .B1(n8030), .C0(n3732), 
        .Y(n3724) );
  INVX3 U8679 ( .A(n3504), .Y(n8456) );
  INVX3 U8680 ( .A(n3299), .Y(n8457) );
  AOI221X2 U8681 ( .A0(n8451), .A1(n7993), .B0(n8452), .B1(n6611), .C0(n3714), 
        .Y(n3706) );
  INVX3 U8682 ( .A(n3503), .Y(n8451) );
  INVX3 U8683 ( .A(n3298), .Y(n8452) );
  AOI221X2 U8684 ( .A0(n8466), .A1(n7993), .B0(n8467), .B1(n6611), .C0(n3750), 
        .Y(n3742) );
  INVX3 U8685 ( .A(n3505), .Y(n8466) );
  INVX3 U8686 ( .A(n3300), .Y(n8467) );
  INVX3 U8687 ( .A(n3500), .Y(n8461) );
  INVX3 U8688 ( .A(n3295), .Y(n8462) );
  AOI2BB2XL U8689 ( .B0(n7982), .B1(n7494), .A0N(n8918), .A1N(n7978), .Y(n3575) );
  AOI2BB2XL U8690 ( .B0(n8047), .B1(n7494), .A0N(n8916), .A1N(n8042), .Y(n3229) );
  AOI2BB2XL U8691 ( .B0(n8098), .B1(n7494), .A0N(n8914), .A1N(n8093), .Y(n2946) );
  AOI2BB2XL U8692 ( .B0(n8111), .B1(n7494), .A0N(n8913), .A1N(n8106), .Y(n2813) );
  AOI2BB2XL U8693 ( .B0(n8123), .B1(n7494), .A0N(n8912), .A1N(n8119), .Y(n2739) );
  AOI2BB2XL U8694 ( .B0(n7969), .B1(n7494), .A0N(n8911), .A1N(n7966), .Y(n3739) );
  AOI2BB2XL U8695 ( .B0(n7982), .B1(n7500), .A0N(n8894), .A1N(n7978), .Y(n3570) );
  AOI2BB2XL U8696 ( .B0(n8046), .B1(n7500), .A0N(n8892), .A1N(n8042), .Y(n3224) );
  AOI2BB2XL U8697 ( .B0(n8098), .B1(n7500), .A0N(n8890), .A1N(n8093), .Y(n2941) );
  AOI2BB2XL U8698 ( .B0(n8111), .B1(n7500), .A0N(n8889), .A1N(n8106), .Y(n2805) );
  AOI2BB2XL U8699 ( .B0(n8123), .B1(n7500), .A0N(n8888), .A1N(n8119), .Y(n2734) );
  AOI2BB2XL U8700 ( .B0(n7969), .B1(n7500), .A0N(n8887), .A1N(n7966), .Y(n3651) );
  AOI2BB2XL U8701 ( .B0(n7982), .B1(n7496), .A0N(n8910), .A1N(n7978), .Y(n3574) );
  AOI2BB2XL U8702 ( .B0(n8046), .B1(n7496), .A0N(n8908), .A1N(n8042), .Y(n3228) );
  AOI2BB2XL U8703 ( .B0(n8098), .B1(n7496), .A0N(n8906), .A1N(n8093), .Y(n2945) );
  AOI2BB2XL U8704 ( .B0(n8111), .B1(n7496), .A0N(n8905), .A1N(n8106), .Y(n2811) );
  AOI2BB2XL U8705 ( .B0(n8123), .B1(n7496), .A0N(n8904), .A1N(n8119), .Y(n2738) );
  AOI2BB2XL U8706 ( .B0(n7970), .B1(n7496), .A0N(n8903), .A1N(n7966), .Y(n3721) );
  AOI2BB2XL U8707 ( .B0(n7982), .B1(n7498), .A0N(n8902), .A1N(n7978), .Y(n3573) );
  AOI2BB2XL U8708 ( .B0(n8046), .B1(n7498), .A0N(n8900), .A1N(n8042), .Y(n3227) );
  AOI2BB2XL U8709 ( .B0(n8098), .B1(n7498), .A0N(n8898), .A1N(n8093), .Y(n2944) );
  AOI2BB2XL U8710 ( .B0(n8111), .B1(n7498), .A0N(n8897), .A1N(n8106), .Y(n2809) );
  AOI2BB2XL U8711 ( .B0(n8123), .B1(n7498), .A0N(n8896), .A1N(n8119), .Y(n2737) );
  AOI2BB2XL U8712 ( .B0(n7969), .B1(n7498), .A0N(n8895), .A1N(n7966), .Y(n3703) );
  NAND2X4 U8713 ( .A(n8885), .B(n8886), .Y(n777) );
  OA22XL U8714 ( .A0(n7760), .A1(n751), .B0(n8350), .B1(n1277), .Y(n1276) );
  OA22X4 U8715 ( .A0(n7758), .A1(n766), .B0(n8347), .B1(n971), .Y(n970) );
  OA22XL U8716 ( .A0(n7754), .A1(n971), .B0(n8340), .B1(n1546), .Y(n1545) );
  INVX3 U8717 ( .A(n2344), .Y(n8469) );
  INVX3 U8718 ( .A(n2534), .Y(n8470) );
  OAI222X2 U8719 ( .A0(n8083), .A1(n3017), .B0(n8019), .B1(n3369), .C0(n8070), 
        .C1(n3088), .Y(n3771) );
  INVX3 U8720 ( .A(n2347), .Y(n8474) );
  INVX3 U8721 ( .A(n2535), .Y(n8475) );
  OAI222X2 U8722 ( .A0(n8083), .A1(n3018), .B0(n8019), .B1(n3370), .C0(n8070), 
        .C1(n3089), .Y(n3789) );
  AOI221X2 U8723 ( .A0(n8471), .A1(n7993), .B0(n8472), .B1(n8030), .C0(n3768), 
        .Y(n3760) );
  INVX3 U8724 ( .A(n3506), .Y(n8471) );
  INVX3 U8725 ( .A(n3301), .Y(n8472) );
  AOI221X2 U8726 ( .A0(n8476), .A1(n6582), .B0(n8477), .B1(n8029), .C0(n3786), 
        .Y(n3778) );
  INVX3 U8727 ( .A(n3507), .Y(n8476) );
  INVX3 U8728 ( .A(n3302), .Y(n8477) );
  AOI2BB2XL U8729 ( .B0(n7982), .B1(n7492), .A0N(n8926), .A1N(n7978), .Y(n3576) );
  AOI2BB2XL U8730 ( .B0(n8048), .B1(n7492), .A0N(n8924), .A1N(n8042), .Y(n3230) );
  AOI2BB2XL U8731 ( .B0(n8098), .B1(n7492), .A0N(n8922), .A1N(n8093), .Y(n2947) );
  AOI2BB2XL U8732 ( .B0(n8111), .B1(n7492), .A0N(n8921), .A1N(n8106), .Y(n2815) );
  AOI2BB2XL U8733 ( .B0(n8123), .B1(n7492), .A0N(n8920), .A1N(n8119), .Y(n2740) );
  AOI2BB2XL U8734 ( .B0(n7970), .B1(n7492), .A0N(n8919), .A1N(n7966), .Y(n3757) );
  AOI2BB2XL U8735 ( .B0(n7982), .B1(n7490), .A0N(n8934), .A1N(n7978), .Y(n3577) );
  AOI2BB2XL U8736 ( .B0(n8045), .B1(n7490), .A0N(n8932), .A1N(n8042), .Y(n3231) );
  AOI2BB2XL U8737 ( .B0(n8098), .B1(n7490), .A0N(n8930), .A1N(n8093), .Y(n2948) );
  AOI2BB2XL U8738 ( .B0(n8111), .B1(n7490), .A0N(n8929), .A1N(n8106), .Y(n2817) );
  AOI2BB2XL U8739 ( .B0(n8123), .B1(n7490), .A0N(n8928), .A1N(n8119), .Y(n2741) );
  AOI2BB2XL U8740 ( .B0(n7970), .B1(n7490), .A0N(n8927), .A1N(n7966), .Y(n3775) );
  OA22XL U8741 ( .A0(n7760), .A1(n743), .B0(n8350), .B1(n1272), .Y(n1271) );
  CLKINVX1 U8742 ( .A(n773), .Y(n8859) );
  OA22XL U8743 ( .A0(n7754), .A1(n974), .B0(n8340), .B1(n1550), .Y(n1549) );
  OA22XL U8744 ( .A0(n7760), .A1(n759), .B0(n8350), .B1(n1282), .Y(n1281) );
  OA22XL U8745 ( .A0(n7753), .A1(n953), .B0(n8341), .B1(n1522), .Y(n1521) );
  OA22XL U8746 ( .A0(n7756), .A1(n1267), .B0(n8345), .B1(n1727), .Y(n1726) );
  OA22XL U8747 ( .A0(n7758), .A1(n734), .B0(n8347), .B1(n959), .Y(n958) );
  INVX3 U8748 ( .A(n2350), .Y(n8479) );
  INVX3 U8749 ( .A(n2536), .Y(n8480) );
  OAI222X2 U8750 ( .A0(n8083), .A1(n3019), .B0(n8019), .B1(n3371), .C0(n8070), 
        .C1(n3090), .Y(n3807) );
  INVX3 U8751 ( .A(n2353), .Y(n8484) );
  INVX3 U8752 ( .A(n2537), .Y(n8485) );
  OAI222X2 U8753 ( .A0(n8083), .A1(n3020), .B0(n8019), .B1(n3372), .C0(n8070), 
        .C1(n3091), .Y(n3825) );
  INVX3 U8754 ( .A(n2356), .Y(n8489) );
  INVX3 U8755 ( .A(n2538), .Y(n8490) );
  OAI222X2 U8756 ( .A0(n8083), .A1(n3021), .B0(n8019), .B1(n3373), .C0(n8070), 
        .C1(n3092), .Y(n3843) );
  AOI221X2 U8757 ( .A0(n8481), .A1(n7994), .B0(n8482), .B1(n8032), .C0(n3804), 
        .Y(n3796) );
  INVX3 U8758 ( .A(n3508), .Y(n8481) );
  INVX3 U8759 ( .A(n3303), .Y(n8482) );
  AOI221X2 U8760 ( .A0(n8486), .A1(n7992), .B0(n8487), .B1(n8032), .C0(n3822), 
        .Y(n3814) );
  INVX3 U8761 ( .A(n3509), .Y(n8486) );
  INVX3 U8762 ( .A(n3304), .Y(n8487) );
  AOI221X2 U8763 ( .A0(n8491), .A1(n7991), .B0(n8492), .B1(n8032), .C0(n3840), 
        .Y(n3832) );
  INVX3 U8764 ( .A(n3510), .Y(n8491) );
  INVX3 U8765 ( .A(n3305), .Y(n8492) );
  AOI2BB2XL U8766 ( .B0(n7982), .B1(n7488), .A0N(n8942), .A1N(n7978), .Y(n3578) );
  AOI2BB2XL U8767 ( .B0(n8046), .B1(n7488), .A0N(n8940), .A1N(n8042), .Y(n3232) );
  AOI2BB2XL U8768 ( .B0(n8098), .B1(n7488), .A0N(n8938), .A1N(n8093), .Y(n2949) );
  AOI2BB2XL U8769 ( .B0(n8111), .B1(n7488), .A0N(n8937), .A1N(n8106), .Y(n2819) );
  AOI2BB2XL U8770 ( .B0(n8123), .B1(n7488), .A0N(n8936), .A1N(n8119), .Y(n2742) );
  AOI2BB2XL U8771 ( .B0(n7969), .B1(n7488), .A0N(n8935), .A1N(n7966), .Y(n3793) );
  AOI2BB2XL U8772 ( .B0(n7982), .B1(n7486), .A0N(n8950), .A1N(n7978), .Y(n3579) );
  AOI2BB2XL U8773 ( .B0(n8046), .B1(n7486), .A0N(n8948), .A1N(n8042), .Y(n3233) );
  AOI2BB2XL U8774 ( .B0(n8098), .B1(n7486), .A0N(n8946), .A1N(n8093), .Y(n2950) );
  AOI2BB2XL U8775 ( .B0(n8111), .B1(n7486), .A0N(n8945), .A1N(n8106), .Y(n2821) );
  AOI2BB2XL U8776 ( .B0(n8123), .B1(n7486), .A0N(n8944), .A1N(n8119), .Y(n2743) );
  AOI2BB2XL U8777 ( .B0(n7970), .B1(n7486), .A0N(n8943), .A1N(n7966), .Y(n3811) );
  AOI2BB2XL U8778 ( .B0(n7982), .B1(n7484), .A0N(n8958), .A1N(n7978), .Y(n3580) );
  AOI2BB2XL U8779 ( .B0(n8046), .B1(n7484), .A0N(n8956), .A1N(n8042), .Y(n3234) );
  AOI2BB2XL U8780 ( .B0(n8098), .B1(n7484), .A0N(n8954), .A1N(n8093), .Y(n2951) );
  AOI2BB2XL U8781 ( .B0(n8111), .B1(n7484), .A0N(n8953), .A1N(n8106), .Y(n2823) );
  AOI2BB2XL U8782 ( .B0(n8123), .B1(n7484), .A0N(n8952), .A1N(n8119), .Y(n2744) );
  AOI2BB2XL U8783 ( .B0(n7969), .B1(n7484), .A0N(n8951), .A1N(n7966), .Y(n3829) );
  OA22XL U8784 ( .A0(n7753), .A1(n947), .B0(n8341), .B1(n1514), .Y(n1513) );
  OA22XL U8785 ( .A0(n7753), .A1(n944), .B0(n8341), .B1(n1510), .Y(n1509) );
  OA22XL U8786 ( .A0(n7755), .A1(n1257), .B0(n8345), .B1(n1721), .Y(n1720) );
  OA22XL U8787 ( .A0(n7755), .A1(n1252), .B0(n8345), .B1(n1718), .Y(n1717) );
  OA22XL U8788 ( .A0(n7757), .A1(n726), .B0(n8347), .B1(n956), .Y(n955) );
  OA22XL U8789 ( .A0(n7757), .A1(n718), .B0(n8347), .B1(n953), .Y(n952) );
  AOI221X2 U8790 ( .A0(n8496), .A1(n7991), .B0(n8497), .B1(n8032), .C0(n3858), 
        .Y(n3850) );
  INVX3 U8791 ( .A(n3511), .Y(n8496) );
  INVX3 U8792 ( .A(n3306), .Y(n8497) );
  AOI221X2 U8793 ( .A0(n8501), .A1(n7991), .B0(n8502), .B1(n8032), .C0(n3876), 
        .Y(n3868) );
  INVX3 U8794 ( .A(n3512), .Y(n8501) );
  INVX3 U8795 ( .A(n3307), .Y(n8502) );
  AOI2BB2XL U8796 ( .B0(n7982), .B1(n7482), .A0N(n8966), .A1N(n7978), .Y(n3581) );
  AOI2BB2XL U8797 ( .B0(n8046), .B1(n7482), .A0N(n8964), .A1N(n8042), .Y(n3235) );
  AOI2BB2XL U8798 ( .B0(n8098), .B1(n7482), .A0N(n8962), .A1N(n8093), .Y(n2952) );
  AOI2BB2XL U8799 ( .B0(n8111), .B1(n7482), .A0N(n8961), .A1N(n8106), .Y(n2825) );
  AOI2BB2XL U8800 ( .B0(n8123), .B1(n7482), .A0N(n8960), .A1N(n8119), .Y(n2745) );
  AOI2BB2XL U8801 ( .B0(n7970), .B1(n7482), .A0N(n8959), .A1N(n7966), .Y(n3847) );
  AOI2BB2XL U8802 ( .B0(n7982), .B1(n7480), .A0N(n8974), .A1N(n7978), .Y(n3582) );
  AOI2BB2XL U8803 ( .B0(n8046), .B1(n7480), .A0N(n8972), .A1N(n8042), .Y(n3236) );
  AOI2BB2XL U8804 ( .B0(n8098), .B1(n7480), .A0N(n8970), .A1N(n8093), .Y(n2953) );
  AOI2BB2XL U8805 ( .B0(n8111), .B1(n7480), .A0N(n8969), .A1N(n8106), .Y(n2827) );
  AOI2BB2XL U8806 ( .B0(n8123), .B1(n7480), .A0N(n8968), .A1N(n8119), .Y(n2746) );
  AOI2BB2XL U8807 ( .B0(n7969), .B1(n7480), .A0N(n8967), .A1N(n7966), .Y(n3865) );
  OA22XL U8808 ( .A0(n7753), .A1(n941), .B0(n8341), .B1(n1506), .Y(n1505) );
  OA22XL U8809 ( .A0(n7759), .A1(n703), .B0(n8350), .B1(n1247), .Y(n1246) );
  OA22XL U8810 ( .A0(n7755), .A1(n1247), .B0(n8345), .B1(n1715), .Y(n1714) );
  OA22XL U8811 ( .A0(n7755), .A1(n1242), .B0(n8345), .B1(n1712), .Y(n1711) );
  OA22XL U8812 ( .A0(n7757), .A1(n710), .B0(n8347), .B1(n950), .Y(n949) );
  AOI221X2 U8813 ( .A0(n8516), .A1(n7991), .B0(n8517), .B1(n8032), .C0(n3930), 
        .Y(n3922) );
  AOI2BB2XL U8814 ( .B0(n7983), .B1(n7474), .A0N(n8998), .A1N(n7979), .Y(n3585) );
  AOI2BB2XL U8815 ( .B0(n8047), .B1(n7474), .A0N(n8996), .A1N(n8043), .Y(n3239) );
  AOI2BB2XL U8816 ( .B0(n8099), .B1(n7474), .A0N(n8994), .A1N(n8094), .Y(n2956) );
  AOI2BB2XL U8817 ( .B0(n8112), .B1(n7474), .A0N(n8993), .A1N(n8107), .Y(n2833) );
  AOI2BB2XL U8818 ( .B0(n8122), .B1(n7474), .A0N(n8992), .A1N(n8120), .Y(n2749) );
  AOI2BB2XL U8819 ( .B0(n7969), .B1(n7474), .A0N(n8991), .A1N(n7967), .Y(n3919) );
  AOI2BB2XL U8820 ( .B0(n7983), .B1(n7472), .A0N(n9006), .A1N(n7979), .Y(n3586) );
  AOI2BB2XL U8821 ( .B0(n8047), .B1(n7472), .A0N(n9004), .A1N(n8043), .Y(n3240) );
  AOI2BB2XL U8822 ( .B0(n8099), .B1(n7472), .A0N(n9002), .A1N(n8094), .Y(n2957) );
  AOI2BB2XL U8823 ( .B0(n8112), .B1(n7472), .A0N(n9001), .A1N(n8107), .Y(n2835) );
  AOI2BB2XL U8824 ( .B0(n8122), .B1(n7472), .A0N(n9000), .A1N(n8120), .Y(n2750) );
  AOI2BB2XL U8825 ( .B0(n7969), .B1(n7472), .A0N(n8999), .A1N(n7967), .Y(n3937) );
  INVXL U8826 ( .A(n3514), .Y(n8511) );
  OA22XL U8827 ( .A0(n7753), .A1(n938), .B0(n8341), .B1(n1502), .Y(n1501) );
  OA22XL U8828 ( .A0(n7759), .A1(n695), .B0(n8350), .B1(n1242), .Y(n1241) );
  OA22XL U8829 ( .A0(n7759), .A1(n687), .B0(n8350), .B1(n1237), .Y(n1236) );
  OA22XL U8830 ( .A0(n7753), .A1(n935), .B0(n8341), .B1(n1498), .Y(n1497) );
  OA22XL U8831 ( .A0(n7755), .A1(n1237), .B0(n8345), .B1(n1709), .Y(n1708) );
  OA22XL U8832 ( .A0(n7757), .A1(n702), .B0(n8347), .B1(n947), .Y(n946) );
  OA22XL U8833 ( .A0(n7757), .A1(n694), .B0(n8347), .B1(n944), .Y(n943) );
  AOI2BB2XL U8834 ( .B0(n7983), .B1(n7470), .A0N(n9014), .A1N(n7979), .Y(n3587) );
  AOI2BB2XL U8835 ( .B0(n8047), .B1(n7470), .A0N(n9012), .A1N(n8043), .Y(n3241) );
  AOI2BB2XL U8836 ( .B0(n8099), .B1(n7470), .A0N(n9010), .A1N(n8094), .Y(n2958) );
  AOI2BB2XL U8837 ( .B0(n8112), .B1(n7470), .A0N(n9009), .A1N(n8107), .Y(n2837) );
  AOI2BB2XL U8838 ( .B0(n8123), .B1(n7470), .A0N(n9008), .A1N(n8120), .Y(n2751) );
  AOI2BB2XL U8839 ( .B0(n7969), .B1(n7470), .A0N(n9007), .A1N(n7967), .Y(n3955) );
  AOI2BB2XL U8840 ( .B0(n7983), .B1(n7468), .A0N(n9022), .A1N(n7979), .Y(n3588) );
  AOI2BB2XL U8841 ( .B0(n8047), .B1(n7468), .A0N(n9020), .A1N(n8043), .Y(n3242) );
  AOI2BB2XL U8842 ( .B0(n8099), .B1(n7468), .A0N(n9018), .A1N(n8094), .Y(n2959) );
  AOI2BB2XL U8843 ( .B0(n8112), .B1(n7468), .A0N(n9017), .A1N(n8107), .Y(n2839) );
  AOI2BB2XL U8844 ( .B0(n8123), .B1(n7468), .A0N(n9016), .A1N(n8120), .Y(n2752) );
  AOI2BB2XL U8845 ( .B0(n7969), .B1(n7468), .A0N(n9015), .A1N(n7967), .Y(n3973) );
  AOI2BB2XL U8846 ( .B0(n7983), .B1(n7466), .A0N(n9030), .A1N(n7979), .Y(n3589) );
  AOI2BB2XL U8847 ( .B0(n8047), .B1(n7466), .A0N(n9028), .A1N(n8043), .Y(n3243) );
  AOI2BB2XL U8848 ( .B0(n8099), .B1(n7466), .A0N(n9026), .A1N(n8094), .Y(n2960) );
  AOI2BB2XL U8849 ( .B0(n8112), .B1(n7466), .A0N(n9025), .A1N(n8107), .Y(n2841) );
  AOI2BB2XL U8850 ( .B0(n8124), .B1(n7466), .A0N(n9024), .A1N(n8120), .Y(n2753) );
  AOI2BB2XL U8851 ( .B0(n7969), .B1(n7466), .A0N(n9023), .A1N(n7967), .Y(n3991) );
  OA22XL U8852 ( .A0(n7759), .A1(n679), .B0(n8350), .B1(n1232), .Y(n1231) );
  OA22XL U8853 ( .A0(n7753), .A1(n932), .B0(n8345), .B1(n1494), .Y(n1493) );
  OA22XL U8854 ( .A0(n7753), .A1(n929), .B0(n8341), .B1(n1490), .Y(n1489) );
  OA22XL U8855 ( .A0(n7759), .A1(n671), .B0(n8350), .B1(n1227), .Y(n1226) );
  OA22XL U8856 ( .A0(n7755), .A1(n1227), .B0(n8345), .B1(n1703), .Y(n1702) );
  OA22XL U8857 ( .A0(n7755), .A1(n1222), .B0(n8345), .B1(n1700), .Y(n1699) );
  OA22XL U8858 ( .A0(n7757), .A1(n686), .B0(n8347), .B1(n941), .Y(n940) );
  OA22XL U8859 ( .A0(n7757), .A1(n678), .B0(n8347), .B1(n938), .Y(n937) );
  INVXL U8860 ( .A(n2392), .Y(n8549) );
  INVXL U8861 ( .A(n2550), .Y(n8550) );
  AOI2BB2XL U8862 ( .B0(n7983), .B1(n7464), .A0N(n9038), .A1N(n7979), .Y(n3590) );
  AOI2BB2XL U8863 ( .B0(n8047), .B1(n7464), .A0N(n9036), .A1N(n8043), .Y(n3244) );
  AOI2BB2XL U8864 ( .B0(n8099), .B1(n7464), .A0N(n9034), .A1N(n8094), .Y(n2961) );
  AOI2BB2XL U8865 ( .B0(n8112), .B1(n7464), .A0N(n9033), .A1N(n8107), .Y(n2843) );
  AOI2BB2XL U8866 ( .B0(n8125), .B1(n7464), .A0N(n9032), .A1N(n8120), .Y(n2754) );
  AOI2BB2XL U8867 ( .B0(n7969), .B1(n7464), .A0N(n9031), .A1N(n7967), .Y(n4009) );
  AOI2BB2XL U8868 ( .B0(n7983), .B1(n7462), .A0N(n9046), .A1N(n7979), .Y(n3591) );
  AOI2BB2XL U8869 ( .B0(n8047), .B1(n7462), .A0N(n9044), .A1N(n8043), .Y(n3245) );
  AOI2BB2XL U8870 ( .B0(n8099), .B1(n7462), .A0N(n9042), .A1N(n8094), .Y(n2962) );
  AOI2BB2XL U8871 ( .B0(n8112), .B1(n7462), .A0N(n9041), .A1N(n8107), .Y(n2845) );
  AOI2BB2XL U8872 ( .B0(n8123), .B1(n7462), .A0N(n9040), .A1N(n8120), .Y(n2755) );
  AOI2BB2XL U8873 ( .B0(n7969), .B1(n7462), .A0N(n9039), .A1N(n7967), .Y(n4027) );
  OA22XL U8874 ( .A0(n7753), .A1(n926), .B0(n8341), .B1(n1486), .Y(n1485) );
  OA22XL U8875 ( .A0(n7759), .A1(n663), .B0(n8350), .B1(n1222), .Y(n1221) );
  OA22XL U8876 ( .A0(n7753), .A1(n923), .B0(n8341), .B1(n1482), .Y(n1481) );
  OA22XL U8877 ( .A0(n7759), .A1(n655), .B0(n8350), .B1(n1217), .Y(n1216) );
  OA22XL U8878 ( .A0(n7757), .A1(n670), .B0(n8347), .B1(n935), .Y(n934) );
  OA22XL U8879 ( .A0(n7755), .A1(n1217), .B0(n8345), .B1(n1697), .Y(n1696) );
  OA22XL U8880 ( .A0(n7757), .A1(n662), .B0(n8347), .B1(n932), .Y(n931) );
  OA22XL U8881 ( .A0(n7755), .A1(n1212), .B0(n8344), .B1(n1694), .Y(n1693) );
  INVXL U8882 ( .A(n2395), .Y(n8554) );
  INVXL U8883 ( .A(n2551), .Y(n8555) );
  INVXL U8884 ( .A(n2398), .Y(n8559) );
  INVXL U8885 ( .A(n2552), .Y(n8560) );
  INVXL U8886 ( .A(n3522), .Y(n8551) );
  INVXL U8887 ( .A(n3317), .Y(n8552) );
  AOI2BB2XL U8888 ( .B0(n7983), .B1(n7457), .A0N(n9070), .A1N(n7979), .Y(n3594) );
  AOI2BB2XL U8889 ( .B0(n8099), .B1(n7457), .A0N(n9066), .A1N(n8094), .Y(n2965) );
  AOI2BB2XL U8890 ( .B0(n8112), .B1(n7457), .A0N(n9065), .A1N(n8107), .Y(n2851) );
  AOI2BB2XL U8891 ( .B0(n8122), .B1(n7457), .A0N(n9064), .A1N(n8120), .Y(n2758) );
  AOI2BB2XL U8892 ( .B0(n7969), .B1(n7457), .A0N(n9063), .A1N(n7967), .Y(n4081) );
  INVXL U8893 ( .A(n3318), .Y(n8557) );
  INVXL U8894 ( .A(n3319), .Y(n8562) );
  INVXL U8895 ( .A(n3523), .Y(n8556) );
  INVXL U8896 ( .A(n3524), .Y(n8561) );
  OA22XL U8897 ( .A0(n7753), .A1(n920), .B0(n8341), .B1(n1478), .Y(n1477) );
  OA22XL U8898 ( .A0(n7759), .A1(n647), .B0(n8350), .B1(n1212), .Y(n1211) );
  OA22XL U8899 ( .A0(n7759), .A1(n639), .B0(n8350), .B1(n1207), .Y(n1206) );
  OA22XL U8900 ( .A0(n7753), .A1(n917), .B0(n8341), .B1(n1474), .Y(n1473) );
  OA22XL U8901 ( .A0(n7757), .A1(n654), .B0(n8347), .B1(n929), .Y(n928) );
  OA22XL U8902 ( .A0(n7755), .A1(n1207), .B0(n8344), .B1(n1691), .Y(n1690) );
  OA22XL U8903 ( .A0(n7757), .A1(n646), .B0(n8346), .B1(n926), .Y(n925) );
  OA22XL U8904 ( .A0(n7755), .A1(n1202), .B0(n8344), .B1(n1688), .Y(n1687) );
  AOI2BB2XL U8905 ( .B0(n7983), .B1(n7455), .A0N(n9078), .A1N(n7979), .Y(n3595) );
  AOI2BB2XL U8906 ( .B0(n8047), .B1(n7455), .A0N(n9076), .A1N(n8043), .Y(n3249) );
  AOI2BB2XL U8907 ( .B0(n8099), .B1(n7455), .A0N(n9074), .A1N(n8094), .Y(n2966) );
  AOI2BB2XL U8908 ( .B0(n8112), .B1(n7455), .A0N(n9073), .A1N(n8107), .Y(n2853) );
  AOI2BB2XL U8909 ( .B0(n8122), .B1(n7455), .A0N(n9072), .A1N(n8120), .Y(n2759) );
  AOI2BB2XL U8910 ( .B0(n7969), .B1(n7455), .A0N(n9071), .A1N(n7967), .Y(n4099) );
  AOI2BB2XL U8911 ( .B0(n7983), .B1(n7453), .A0N(n9086), .A1N(n7980), .Y(n3596) );
  AOI2BB2XL U8912 ( .B0(n8047), .B1(n7453), .A0N(n9084), .A1N(n8044), .Y(n3250) );
  AOI2BB2XL U8913 ( .B0(n8099), .B1(n7453), .A0N(n9082), .A1N(n8095), .Y(n2967) );
  AOI2BB2XL U8914 ( .B0(n8112), .B1(n7453), .A0N(n9081), .A1N(n8108), .Y(n2855) );
  AOI2BB2XL U8915 ( .B0(n8122), .B1(n7453), .A0N(n9080), .A1N(n8121), .Y(n2760) );
  AOI2BB2XL U8916 ( .B0(n7969), .B1(n7453), .A0N(n9079), .A1N(n7968), .Y(n4117) );
  AOI2BB2XL U8917 ( .B0(n7983), .B1(n7451), .A0N(n9094), .A1N(n7980), .Y(n3597) );
  AOI2BB2XL U8918 ( .B0(n8047), .B1(n7451), .A0N(n9092), .A1N(n8044), .Y(n3251) );
  AOI2BB2XL U8919 ( .B0(n8099), .B1(n7451), .A0N(n9090), .A1N(n8095), .Y(n2968) );
  AOI2BB2XL U8920 ( .B0(n8112), .B1(n7451), .A0N(n9089), .A1N(n8108), .Y(n2857) );
  AOI2BB2XL U8921 ( .B0(n8122), .B1(n7451), .A0N(n9088), .A1N(n8121), .Y(n2761) );
  AOI2BB2XL U8922 ( .B0(n7969), .B1(n7451), .A0N(n9087), .A1N(n7968), .Y(n4135) );
  OA22XL U8923 ( .A0(n7753), .A1(n911), .B0(n8341), .B1(n1466), .Y(n1465) );
  OA22XL U8924 ( .A0(n7753), .A1(n914), .B0(n8341), .B1(n1470), .Y(n1469) );
  OA22XL U8925 ( .A0(n7759), .A1(n631), .B0(n8349), .B1(n1202), .Y(n1201) );
  OA22XL U8926 ( .A0(n7759), .A1(n623), .B0(n8349), .B1(n1197), .Y(n1196) );
  OA22XL U8927 ( .A0(n7755), .A1(n1197), .B0(n8344), .B1(n1685), .Y(n1684) );
  OA22XL U8928 ( .A0(n7757), .A1(n630), .B0(n8346), .B1(n920), .Y(n919) );
  OA22XL U8929 ( .A0(n7755), .A1(n1192), .B0(n8344), .B1(n1682), .Y(n1681) );
  AOI2BB2XL U8930 ( .B0(n7984), .B1(n7449), .A0N(n9102), .A1N(n7980), .Y(n3598) );
  AOI2BB2XL U8931 ( .B0(n8048), .B1(n7449), .A0N(n9100), .A1N(n8044), .Y(n3252) );
  AOI2BB2XL U8932 ( .B0(n8096), .B1(n7449), .A0N(n9098), .A1N(n8095), .Y(n2969) );
  AOI2BB2XL U8933 ( .B0(n8110), .B1(n7449), .A0N(n9097), .A1N(n8108), .Y(n2859) );
  AOI2BB2XL U8934 ( .B0(n8124), .B1(n7449), .A0N(n9096), .A1N(n8121), .Y(n2762) );
  AOI2BB2XL U8935 ( .B0(n7970), .B1(n7449), .A0N(n9095), .A1N(n7968), .Y(n4153) );
  AOI2BB2XL U8936 ( .B0(n7984), .B1(n7447), .A0N(n9110), .A1N(n7980), .Y(n3599) );
  AOI2BB2XL U8937 ( .B0(n8048), .B1(n7447), .A0N(n9108), .A1N(n8044), .Y(n3253) );
  AOI2BB2XL U8938 ( .B0(n8096), .B1(n7447), .A0N(n9106), .A1N(n8095), .Y(n2970) );
  AOI2BB2XL U8939 ( .B0(n8110), .B1(n7447), .A0N(n9105), .A1N(n8108), .Y(n2861) );
  AOI2BB2XL U8940 ( .B0(n8124), .B1(n7447), .A0N(n9104), .A1N(n8121), .Y(n2763) );
  AOI2BB2XL U8941 ( .B0(n7970), .B1(n7447), .A0N(n9103), .A1N(n7968), .Y(n4171) );
  AOI2BB2XL U8942 ( .B0(n7984), .B1(n7445), .A0N(n9118), .A1N(n7980), .Y(n3600) );
  AOI2BB2XL U8943 ( .B0(n8048), .B1(n7445), .A0N(n9116), .A1N(n8044), .Y(n3254) );
  AOI2BB2XL U8944 ( .B0(n8096), .B1(n7445), .A0N(n9114), .A1N(n8095), .Y(n2971) );
  AOI2BB2XL U8945 ( .B0(n8110), .B1(n7445), .A0N(n9113), .A1N(n8108), .Y(n2863) );
  AOI2BB2XL U8946 ( .B0(n8124), .B1(n7445), .A0N(n9112), .A1N(n8121), .Y(n2764) );
  AOI2BB2XL U8947 ( .B0(n7970), .B1(n7445), .A0N(n9111), .A1N(n7968), .Y(n4189) );
  OA22XL U8948 ( .A0(n7753), .A1(n905), .B0(n8341), .B1(n1458), .Y(n1457) );
  OA22XL U8949 ( .A0(n7753), .A1(n908), .B0(n8341), .B1(n1462), .Y(n1461) );
  OA22XL U8950 ( .A0(n7759), .A1(n607), .B0(n8349), .B1(n1187), .Y(n1186) );
  OA22XL U8951 ( .A0(n7759), .A1(n615), .B0(n8349), .B1(n1192), .Y(n1191) );
  OA22XL U8952 ( .A0(n7757), .A1(n622), .B0(n8346), .B1(n917), .Y(n916) );
  OA22XL U8953 ( .A0(n7755), .A1(n1187), .B0(n8344), .B1(n1679), .Y(n1678) );
  OA22XL U8954 ( .A0(n7757), .A1(n614), .B0(n8346), .B1(n914), .Y(n913) );
  INVXL U8955 ( .A(n2425), .Y(n8604) );
  INVXL U8956 ( .A(n2561), .Y(n8605) );
  AOI2BB2XL U8957 ( .B0(n7984), .B1(n7443), .A0N(n9126), .A1N(n7980), .Y(n3601) );
  AOI2BB2XL U8958 ( .B0(n8048), .B1(n7443), .A0N(n9124), .A1N(n8044), .Y(n3255) );
  AOI2BB2XL U8959 ( .B0(n8096), .B1(n7443), .A0N(n9122), .A1N(n8095), .Y(n2972) );
  AOI2BB2XL U8960 ( .B0(n8110), .B1(n7443), .A0N(n9121), .A1N(n8108), .Y(n2865) );
  AOI2BB2XL U8961 ( .B0(n8124), .B1(n7443), .A0N(n9120), .A1N(n8121), .Y(n2765) );
  AOI2BB2XL U8962 ( .B0(n7970), .B1(n7443), .A0N(n9119), .A1N(n7968), .Y(n4207) );
  AOI2BB2XL U8963 ( .B0(n7984), .B1(n7441), .A0N(n9134), .A1N(n7980), .Y(n3602) );
  AOI2BB2XL U8964 ( .B0(n8048), .B1(n7441), .A0N(n9132), .A1N(n8044), .Y(n3256) );
  AOI2BB2XL U8965 ( .B0(n8096), .B1(n7441), .A0N(n9130), .A1N(n8095), .Y(n2973) );
  AOI2BB2XL U8966 ( .B0(n8109), .B1(n7441), .A0N(n9129), .A1N(n8108), .Y(n2867) );
  AOI2BB2XL U8967 ( .B0(n8124), .B1(n7441), .A0N(n9128), .A1N(n8121), .Y(n2766) );
  AOI2BB2XL U8968 ( .B0(n7970), .B1(n7441), .A0N(n9127), .A1N(n7968), .Y(n4225) );
  AOI2BB2XL U8969 ( .B0(n7984), .B1(n7439), .A0N(n9142), .A1N(n7980), .Y(n3603) );
  AOI2BB2XL U8970 ( .B0(n8099), .B1(n7439), .A0N(n9138), .A1N(n8095), .Y(n2974) );
  AOI2BB2XL U8971 ( .B0(n8110), .B1(n7439), .A0N(n9137), .A1N(n8108), .Y(n2869) );
  AOI2BB2XL U8972 ( .B0(n8124), .B1(n7439), .A0N(n9136), .A1N(n8121), .Y(n2767) );
  AOI2BB2XL U8973 ( .B0(n7970), .B1(n7439), .A0N(n9135), .A1N(n7968), .Y(n4243) );
  INVXL U8974 ( .A(n3328), .Y(n8607) );
  OA22XL U8975 ( .A0(n7752), .A1(n899), .B0(n8341), .B1(n1450), .Y(n1449) );
  OA22XL U8976 ( .A0(n7753), .A1(n902), .B0(n8341), .B1(n1454), .Y(n1453) );
  OA22XL U8977 ( .A0(n7759), .A1(n591), .B0(n8349), .B1(n1177), .Y(n1176) );
  OA22XL U8978 ( .A0(n7759), .A1(n599), .B0(n8349), .B1(n1182), .Y(n1181) );
  OA22XL U8979 ( .A0(n7757), .A1(n606), .B0(n8346), .B1(n911), .Y(n910) );
  OA22XL U8980 ( .A0(n7755), .A1(n1177), .B0(n8344), .B1(n1673), .Y(n1672) );
  OA22XL U8981 ( .A0(n7757), .A1(n598), .B0(n8346), .B1(n908), .Y(n907) );
  INVXL U8982 ( .A(n2428), .Y(n8609) );
  INVXL U8983 ( .A(n2562), .Y(n8610) );
  AOI2BB2XL U8984 ( .B0(n8124), .B1(n7437), .A0N(n9144), .A1N(n8121), .Y(n2768) );
  AOI2BB2XL U8985 ( .B0(n7984), .B1(n7435), .A0N(n9158), .A1N(n7980), .Y(n3605) );
  AOI2BB2XL U8986 ( .B0(n8048), .B1(n7435), .A0N(n9156), .A1N(n8044), .Y(n3259) );
  AOI2BB2XL U8987 ( .B0(n8096), .B1(n7435), .A0N(n9154), .A1N(n8095), .Y(n2976) );
  AOI2BB2XL U8988 ( .B0(n8110), .B1(n7435), .A0N(n9153), .A1N(n8108), .Y(n2873) );
  AOI2BB2XL U8989 ( .B0(n8124), .B1(n7435), .A0N(n9152), .A1N(n8121), .Y(n2769) );
  AOI2BB2XL U8990 ( .B0(n7970), .B1(n7435), .A0N(n9151), .A1N(n7968), .Y(n4279) );
  AOI2BB2XL U8991 ( .B0(n7984), .B1(n7433), .A0N(n9166), .A1N(n7980), .Y(n3606) );
  AOI2BB2XL U8992 ( .B0(n8048), .B1(n7433), .A0N(n9164), .A1N(n8044), .Y(n3260) );
  AOI2BB2XL U8993 ( .B0(n8096), .B1(n7433), .A0N(n9162), .A1N(n8095), .Y(n2977) );
  AOI2BB2XL U8994 ( .B0(n8110), .B1(n7433), .A0N(n9161), .A1N(n8108), .Y(n2875) );
  AOI2BB2XL U8995 ( .B0(n8124), .B1(n7433), .A0N(n9160), .A1N(n8121), .Y(n2770) );
  AOI2BB2XL U8996 ( .B0(n7970), .B1(n7433), .A0N(n9159), .A1N(n7968), .Y(n4297) );
  INVXL U8997 ( .A(n3329), .Y(n8612) );
  INVXL U8998 ( .A(n3533), .Y(n8606) );
  INVXL U8999 ( .A(n3534), .Y(n8611) );
  OA22XL U9000 ( .A0(n7752), .A1(n893), .B0(n8342), .B1(n1442), .Y(n1441) );
  OA22XL U9001 ( .A0(n7752), .A1(n896), .B0(n8341), .B1(n1446), .Y(n1445) );
  OA22XL U9002 ( .A0(n7759), .A1(n575), .B0(n8349), .B1(n1167), .Y(n1166) );
  OA22XL U9003 ( .A0(n7759), .A1(n583), .B0(n8349), .B1(n1172), .Y(n1171) );
  OA22XL U9004 ( .A0(n7755), .A1(n1172), .B0(n8344), .B1(n1670), .Y(n1669) );
  OA22XL U9005 ( .A0(n7757), .A1(n590), .B0(n8346), .B1(n905), .Y(n904) );
  OA22XL U9006 ( .A0(n7755), .A1(n1167), .B0(n8344), .B1(n1667), .Y(n1666) );
  OA22XL U9007 ( .A0(n7757), .A1(n582), .B0(n8346), .B1(n902), .Y(n901) );
  AOI2BB2XL U9008 ( .B0(n7984), .B1(n7431), .A0N(n9174), .A1N(n7980), .Y(n3607) );
  AOI2BB2XL U9009 ( .B0(n8048), .B1(n7431), .A0N(n9172), .A1N(n8044), .Y(n3261) );
  AOI2BB2XL U9010 ( .B0(n8096), .B1(n7431), .A0N(n9170), .A1N(n8095), .Y(n2978) );
  AOI2BB2XL U9011 ( .B0(n8111), .B1(n7431), .A0N(n9169), .A1N(n8108), .Y(n2877) );
  AOI2BB2XL U9012 ( .B0(n8124), .B1(n7431), .A0N(n9168), .A1N(n8121), .Y(n2771) );
  AOI2BB2XL U9013 ( .B0(n7970), .B1(n7431), .A0N(n9167), .A1N(n7968), .Y(n4315) );
  AOI2BB2XL U9014 ( .B0(n7984), .B1(n7429), .A0N(n9182), .A1N(n7980), .Y(n3608) );
  AOI2BB2XL U9015 ( .B0(n8048), .B1(n7429), .A0N(n9180), .A1N(n8043), .Y(n3262) );
  AOI2BB2XL U9016 ( .B0(n8096), .B1(n7429), .A0N(n9178), .A1N(n8093), .Y(n2979) );
  AOI2BB2XL U9017 ( .B0(n8110), .B1(n7429), .A0N(n9177), .A1N(n8107), .Y(n2879) );
  AOI2BB2XL U9018 ( .B0(n8124), .B1(n7429), .A0N(n9176), .A1N(n8119), .Y(n2772) );
  AOI2BB2XL U9019 ( .B0(n7970), .B1(n7429), .A0N(n9175), .A1N(n7968), .Y(n4333) );
  OA22XL U9020 ( .A0(n7752), .A1(n890), .B0(n8342), .B1(n1438), .Y(n1437) );
  OA22XL U9021 ( .A0(n7759), .A1(n559), .B0(n8349), .B1(n1157), .Y(n1156) );
  OA22XL U9022 ( .A0(n7759), .A1(n567), .B0(n8349), .B1(n1162), .Y(n1161) );
  OA22XL U9023 ( .A0(n7757), .A1(n566), .B0(n8346), .B1(n896), .Y(n895) );
  OA22XL U9024 ( .A0(n7757), .A1(n574), .B0(n8346), .B1(n899), .Y(n898) );
  OA22XL U9025 ( .A0(n7755), .A1(n1162), .B0(n8344), .B1(n1664), .Y(n1663) );
  OA22XL U9026 ( .A0(n7744), .A1(n1157), .B0(n8344), .B1(n1661), .Y(n1660) );
  AOI2BB2XL U9027 ( .B0(n7984), .B1(n7427), .A0N(n9190), .A1N(n7980), .Y(n3609) );
  AOI2BB2XL U9028 ( .B0(n8048), .B1(n7427), .A0N(n9188), .A1N(n8042), .Y(n3263) );
  AOI2BB2XL U9029 ( .B0(n8096), .B1(n7427), .A0N(n9186), .A1N(n8094), .Y(n2980) );
  AOI2BB2XL U9030 ( .B0(n8110), .B1(n7427), .A0N(n9185), .A1N(n2808), .Y(n2881) );
  AOI2BB2XL U9031 ( .B0(n8124), .B1(n7427), .A0N(n9184), .A1N(n8121), .Y(n2773) );
  AOI2BB2XL U9032 ( .B0(n7970), .B1(n7427), .A0N(n9183), .A1N(n7966), .Y(n4351) );
  AOI2BB2XL U9033 ( .B0(n7984), .B1(n7425), .A0N(n9198), .A1N(n7978), .Y(n3610) );
  AOI2BB2XL U9034 ( .B0(n8048), .B1(n7425), .A0N(n9196), .A1N(n8044), .Y(n3264) );
  AOI2BB2XL U9035 ( .B0(n8098), .B1(n7425), .A0N(n9194), .A1N(n8095), .Y(n2981) );
  AOI2BB2XL U9036 ( .B0(n8112), .B1(n7425), .A0N(n9193), .A1N(n8106), .Y(n2883) );
  AOI2BB2XL U9037 ( .B0(n8124), .B1(n7425), .A0N(n9192), .A1N(n8120), .Y(n2774) );
  AOI2BB2XL U9038 ( .B0(n7970), .B1(n7425), .A0N(n9191), .A1N(n7967), .Y(n4369) );
  AOI2BB2XL U9039 ( .B0(n7982), .B1(n7423), .A0N(n9206), .A1N(n7979), .Y(n3611) );
  AOI2BB2XL U9040 ( .B0(n8047), .B1(n7423), .A0N(n9204), .A1N(n8043), .Y(n3265) );
  AOI2BB2XL U9041 ( .B0(n8099), .B1(n7423), .A0N(n9202), .A1N(n8093), .Y(n2982) );
  AOI2BB2XL U9042 ( .B0(n8109), .B1(n7423), .A0N(n9201), .A1N(n8108), .Y(n2885) );
  AOI2BB2XL U9043 ( .B0(n8125), .B1(n7423), .A0N(n9200), .A1N(n8121), .Y(n2775) );
  AOI2BB2XL U9044 ( .B0(n7971), .B1(n7423), .A0N(n9199), .A1N(n7968), .Y(n4387) );
  OA22XL U9045 ( .A0(n7752), .A1(n887), .B0(n8342), .B1(n1434), .Y(n1433) );
  OA22XL U9046 ( .A0(n7752), .A1(n884), .B0(n8342), .B1(n1430), .Y(n1429) );
  OA22XL U9047 ( .A0(n7746), .A1(n551), .B0(n8349), .B1(n1152), .Y(n1151) );
  OA22XL U9048 ( .A0(n7745), .A1(n1147), .B0(n8344), .B1(n1655), .Y(n1654) );
  OA22XL U9049 ( .A0(n7745), .A1(n1152), .B0(n8344), .B1(n1658), .Y(n1657) );
  AOI2BB2XL U9050 ( .B0(n7983), .B1(n7421), .A0N(n9214), .A1N(n3572), .Y(n3612) );
  AOI2BB2XL U9051 ( .B0(n8045), .B1(n7421), .A0N(n9212), .A1N(n3226), .Y(n3266) );
  AOI2BB2XL U9052 ( .B0(n8098), .B1(n7421), .A0N(n9210), .A1N(n8094), .Y(n2983) );
  AOI2BB2XL U9053 ( .B0(n8109), .B1(n7421), .A0N(n9209), .A1N(n8107), .Y(n2887) );
  AOI2BB2XL U9054 ( .B0(n8125), .B1(n7421), .A0N(n9208), .A1N(n8119), .Y(n2776) );
  AOI2BB2XL U9055 ( .B0(n7971), .B1(n7421), .A0N(n9207), .A1N(n7966), .Y(n4405) );
  AOI2BB2XL U9056 ( .B0(n7981), .B1(n7419), .A0N(n9222), .A1N(n7980), .Y(n3613) );
  AOI2BB2XL U9057 ( .B0(n8045), .B1(n7419), .A0N(n9220), .A1N(n8042), .Y(n3267) );
  AOI2BB2XL U9058 ( .B0(n8096), .B1(n7419), .A0N(n9218), .A1N(n8095), .Y(n2984) );
  AOI2BB2XL U9059 ( .B0(n8109), .B1(n7419), .A0N(n9217), .A1N(n8106), .Y(n2889) );
  AOI2BB2XL U9060 ( .B0(n8125), .B1(n7419), .A0N(n9216), .A1N(n8121), .Y(n2777) );
  AOI2BB2XL U9061 ( .B0(n7971), .B1(n7419), .A0N(n9215), .A1N(n7967), .Y(n4423) );
  AOI2BB2XL U9062 ( .B0(n7984), .B1(n7417), .A0N(n9230), .A1N(n7979), .Y(n3614) );
  AOI2BB2XL U9063 ( .B0(n8045), .B1(n7417), .A0N(n9228), .A1N(n8044), .Y(n3268) );
  AOI2BB2XL U9064 ( .B0(n8097), .B1(n7417), .A0N(n9226), .A1N(n2943), .Y(n2985) );
  AOI2BB2XL U9065 ( .B0(n8109), .B1(n7417), .A0N(n9225), .A1N(n2808), .Y(n2891) );
  AOI2BB2XL U9066 ( .B0(n8125), .B1(n7417), .A0N(n9224), .A1N(n8120), .Y(n2778) );
  AOI2BB2XL U9067 ( .B0(n7971), .B1(n7417), .A0N(n9223), .A1N(n3654), .Y(n4441) );
  OA22XL U9068 ( .A0(n7751), .A1(n543), .B0(n8349), .B1(n1147), .Y(n1146) );
  OA22XL U9069 ( .A0(n7741), .A1(n535), .B0(n8349), .B1(n1142), .Y(n1141) );
  OA22XL U9070 ( .A0(n7746), .A1(n881), .B0(n8342), .B1(n1426), .Y(n1425) );
  OA22XL U9071 ( .A0(n7744), .A1(n878), .B0(n8342), .B1(n1422), .Y(n1421) );
  OA22XL U9072 ( .A0(n7745), .A1(n1137), .B0(n8344), .B1(n1649), .Y(n1648) );
  OA22XL U9073 ( .A0(n7750), .A1(n542), .B0(n8346), .B1(n887), .Y(n886) );
  OA22XL U9074 ( .A0(n7745), .A1(n1142), .B0(n8344), .B1(n1652), .Y(n1651) );
  OA22XL U9075 ( .A0(n7751), .A1(n550), .B0(n8346), .B1(n890), .Y(n889) );
  AOI2BB2XL U9076 ( .B0(n7981), .B1(n7415), .A0N(n9238), .A1N(n7978), .Y(n3615) );
  AOI2BB2XL U9077 ( .B0(n8045), .B1(n7415), .A0N(n9236), .A1N(n8043), .Y(n3269) );
  AOI2BB2XL U9078 ( .B0(n8097), .B1(n7415), .A0N(n9234), .A1N(n8095), .Y(n2986) );
  AOI2BB2XL U9079 ( .B0(n8109), .B1(n7415), .A0N(n9233), .A1N(n8108), .Y(n2893) );
  AOI2BB2XL U9080 ( .B0(n8125), .B1(n7415), .A0N(n9232), .A1N(n8120), .Y(n2779) );
  AOI2BB2XL U9081 ( .B0(n7971), .B1(n7415), .A0N(n9231), .A1N(n7966), .Y(n4459) );
  AOI2BB2XL U9082 ( .B0(n7981), .B1(n7413), .A0N(n9246), .A1N(n7979), .Y(n3616) );
  AOI2BB2XL U9083 ( .B0(n8045), .B1(n7413), .A0N(n9244), .A1N(n8043), .Y(n3270) );
  AOI2BB2XL U9084 ( .B0(n8097), .B1(n7413), .A0N(n9242), .A1N(n8095), .Y(n2987) );
  AOI2BB2XL U9085 ( .B0(n8109), .B1(n7413), .A0N(n9241), .A1N(n8107), .Y(n2895) );
  AOI2BB2XL U9086 ( .B0(n8125), .B1(n7413), .A0N(n9240), .A1N(n8121), .Y(n2780) );
  AOI2BB2XL U9087 ( .B0(n7971), .B1(n7413), .A0N(n9239), .A1N(n7968), .Y(n4477) );
  AOI2BB2XL U9088 ( .B0(n7981), .B1(n7411), .A0N(n9254), .A1N(n7980), .Y(n3617) );
  AOI2BB2XL U9089 ( .B0(n8045), .B1(n7411), .A0N(n9252), .A1N(n8042), .Y(n3271) );
  AOI2BB2XL U9090 ( .B0(n8097), .B1(n7411), .A0N(n9250), .A1N(n8093), .Y(n2988) );
  AOI2BB2XL U9091 ( .B0(n8109), .B1(n7411), .A0N(n9249), .A1N(n8107), .Y(n2897) );
  AOI2BB2XL U9092 ( .B0(n8125), .B1(n7411), .A0N(n9248), .A1N(n8119), .Y(n2781) );
  AOI2BB2XL U9093 ( .B0(n7971), .B1(n7411), .A0N(n9247), .A1N(n7966), .Y(n4495) );
  CLKBUFX2 U9094 ( .A(n8410), .Y(n7211) );
  OA22XL U9095 ( .A0(n7741), .A1(n527), .B0(n8349), .B1(n1137), .Y(n1136) );
  OA22XL U9096 ( .A0(n7741), .A1(n519), .B0(n8349), .B1(n1132), .Y(n1131) );
  OA22XL U9097 ( .A0(n7751), .A1(n875), .B0(n8342), .B1(n1418), .Y(n1417) );
  OA22XL U9098 ( .A0(n7746), .A1(n872), .B0(n8342), .B1(n1414), .Y(n1413) );
  OA22XL U9099 ( .A0(n7745), .A1(n1127), .B0(n8344), .B1(n1643), .Y(n1642) );
  OA22XL U9100 ( .A0(n7744), .A1(n526), .B0(n8346), .B1(n881), .Y(n880) );
  OA22XL U9101 ( .A0(n7750), .A1(n534), .B0(n8346), .B1(n884), .Y(n883) );
  AOI2BB2XL U9102 ( .B0(n7981), .B1(n7409), .A0N(n9262), .A1N(n7978), .Y(n3618) );
  AOI2BB2XL U9103 ( .B0(n8045), .B1(n7409), .A0N(n9260), .A1N(n8042), .Y(n3272) );
  AOI2BB2XL U9104 ( .B0(n8097), .B1(n7409), .A0N(n9258), .A1N(n8094), .Y(n2989) );
  AOI2BB2XL U9105 ( .B0(n8109), .B1(n7409), .A0N(n9257), .A1N(n8106), .Y(n2899) );
  AOI2BB2XL U9106 ( .B0(n8125), .B1(n7409), .A0N(n9256), .A1N(n8120), .Y(n2782) );
  AOI2BB2XL U9107 ( .B0(n7971), .B1(n7409), .A0N(n9255), .A1N(n7967), .Y(n4513) );
  AOI2BB2XL U9108 ( .B0(n7981), .B1(n7407), .A0N(n9270), .A1N(n7979), .Y(n3619) );
  AOI2BB2XL U9109 ( .B0(n8045), .B1(n7407), .A0N(n9268), .A1N(n8044), .Y(n3273) );
  AOI2BB2XL U9110 ( .B0(n8097), .B1(n7407), .A0N(n9266), .A1N(n8095), .Y(n2990) );
  AOI2BB2XL U9111 ( .B0(n8109), .B1(n7407), .A0N(n9265), .A1N(n8108), .Y(n2901) );
  AOI2BB2XL U9112 ( .B0(n8125), .B1(n7407), .A0N(n9264), .A1N(n2736), .Y(n2783) );
  AOI2BB2XL U9113 ( .B0(n7969), .B1(n7407), .A0N(n9263), .A1N(n3654), .Y(n4531) );
  AOI2BB2XL U9114 ( .B0(n7981), .B1(n7405), .A0N(n9278), .A1N(n7980), .Y(n3620) );
  AOI2BB2XL U9115 ( .B0(n8045), .B1(n7405), .A0N(n9276), .A1N(n8044), .Y(n3274) );
  AOI2BB2XL U9116 ( .B0(n8097), .B1(n7405), .A0N(n9274), .A1N(n8093), .Y(n2991) );
  AOI2BB2XL U9117 ( .B0(n8109), .B1(n7405), .A0N(n9273), .A1N(n8108), .Y(n2903) );
  AOI2BB2XL U9118 ( .B0(n8125), .B1(n7405), .A0N(n9272), .A1N(n8120), .Y(n2784) );
  AOI2BB2XL U9119 ( .B0(n7970), .B1(n7405), .A0N(n9271), .A1N(n7967), .Y(n4549) );
  OA22XL U9120 ( .A0(n7741), .A1(n511), .B0(n8349), .B1(n1127), .Y(n1126) );
  OA22XL U9121 ( .A0(n7741), .A1(n503), .B0(n8349), .B1(n1122), .Y(n1121) );
  OA22XL U9122 ( .A0(n7744), .A1(n866), .B0(n8342), .B1(n1406), .Y(n1405) );
  OA22XL U9123 ( .A0(n7750), .A1(n869), .B0(n8342), .B1(n1410), .Y(n1409) );
  OA22XL U9124 ( .A0(n7745), .A1(n1117), .B0(n8344), .B1(n1637), .Y(n1636) );
  OA22XL U9125 ( .A0(n7750), .A1(n510), .B0(n8346), .B1(n875), .Y(n874) );
  OA22XL U9126 ( .A0(n7745), .A1(n1122), .B0(n8344), .B1(n1640), .Y(n1639) );
  OA22XL U9127 ( .A0(n7746), .A1(n518), .B0(n8346), .B1(n878), .Y(n877) );
  AOI2BB2XL U9128 ( .B0(n7983), .B1(n7403), .A0N(n9286), .A1N(n7979), .Y(n3621) );
  AOI2BB2XL U9129 ( .B0(n8045), .B1(n7403), .A0N(n9284), .A1N(n8043), .Y(n3275) );
  AOI2BB2XL U9130 ( .B0(n8097), .B1(n7403), .A0N(n9282), .A1N(n8094), .Y(n2992) );
  AOI2BB2XL U9131 ( .B0(n8109), .B1(n7403), .A0N(n9281), .A1N(n8106), .Y(n2905) );
  AOI2BB2XL U9132 ( .B0(n8125), .B1(n7403), .A0N(n9280), .A1N(n2736), .Y(n2785) );
  AOI2BB2XL U9133 ( .B0(n3652), .B1(n7403), .A0N(n9279), .A1N(n7968), .Y(n4567) );
  AOI2BB2XL U9134 ( .B0(n7982), .B1(n7401), .A0N(n9294), .A1N(n7980), .Y(n3622) );
  AOI2BB2XL U9135 ( .B0(n8045), .B1(n7401), .A0N(n9292), .A1N(n8042), .Y(n3276) );
  AOI2BB2XL U9136 ( .B0(n8097), .B1(n7401), .A0N(n9290), .A1N(n8095), .Y(n2993) );
  AOI2BB2XL U9137 ( .B0(n8109), .B1(n7401), .A0N(n9289), .A1N(n8107), .Y(n2907) );
  AOI2BB2XL U9138 ( .B0(n8125), .B1(n7401), .A0N(n9288), .A1N(n2736), .Y(n2786) );
  AOI2BB2XL U9139 ( .B0(n3652), .B1(n7401), .A0N(n9287), .A1N(n7966), .Y(n4585) );
  OA22XL U9140 ( .A0(n7741), .A1(n495), .B0(n8349), .B1(n1117), .Y(n1116) );
  OA22XL U9141 ( .A0(n7741), .A1(n487), .B0(n8349), .B1(n1112), .Y(n1111) );
  OA22XL U9142 ( .A0(n7746), .A1(n860), .B0(n8342), .B1(n1398), .Y(n1397) );
  OA22XL U9143 ( .A0(n7750), .A1(n863), .B0(n8342), .B1(n1402), .Y(n1401) );
  OA22XL U9144 ( .A0(n7745), .A1(n1107), .B0(n8343), .B1(n1631), .Y(n1630) );
  OA22XL U9145 ( .A0(n7750), .A1(n494), .B0(n8346), .B1(n869), .Y(n868) );
  OA22XL U9146 ( .A0(n7745), .A1(n1112), .B0(n8344), .B1(n1634), .Y(n1633) );
  OA22XL U9147 ( .A0(n7744), .A1(n502), .B0(n8346), .B1(n872), .Y(n871) );
  AOI2BB2XL U9148 ( .B0(n7984), .B1(n7399), .A0N(n9302), .A1N(n7978), .Y(n3623) );
  AOI2BB2XL U9149 ( .B0(n8045), .B1(n7399), .A0N(n9300), .A1N(n8044), .Y(n3277) );
  AOI2BB2XL U9150 ( .B0(n8097), .B1(n7399), .A0N(n9298), .A1N(n8093), .Y(n2994) );
  AOI2BB2XL U9151 ( .B0(n8109), .B1(n7399), .A0N(n9297), .A1N(n8108), .Y(n2909) );
  AOI2BB2XL U9152 ( .B0(n8125), .B1(n7399), .A0N(n9296), .A1N(n2736), .Y(n2787) );
  AOI2BB2XL U9153 ( .B0(n7970), .B1(n7399), .A0N(n9295), .A1N(n7968), .Y(n4603) );
  AOI2BB2XL U9154 ( .B0(n3571), .B1(n7397), .A0N(n9310), .A1N(n7978), .Y(n3624) );
  AOI2BB2XL U9155 ( .B0(n3225), .B1(n7397), .A0N(n9308), .A1N(n8042), .Y(n3278) );
  AOI2BB2XL U9156 ( .B0(n2942), .B1(n7397), .A0N(n9306), .A1N(n8093), .Y(n2995) );
  AOI2BB2XL U9157 ( .B0(n2806), .B1(n7397), .A0N(n9305), .A1N(n8108), .Y(n2911) );
  AOI2BB2XL U9158 ( .B0(n8122), .B1(n7397), .A0N(n9304), .A1N(n8121), .Y(n2788) );
  AOI2BB2XL U9159 ( .B0(n7971), .B1(n7397), .A0N(n9303), .A1N(n7967), .Y(n4621) );
  AOI2BB2XL U9160 ( .B0(n7981), .B1(n7395), .A0N(n9318), .A1N(n7978), .Y(n3625) );
  AOI2BB2XL U9161 ( .B0(n8046), .B1(n7395), .A0N(n9316), .A1N(n8043), .Y(n3279) );
  AOI2BB2XL U9162 ( .B0(n2942), .B1(n7395), .A0N(n9314), .A1N(n8094), .Y(n2996) );
  AOI2BB2XL U9163 ( .B0(n8110), .B1(n7395), .A0N(n9313), .A1N(n8106), .Y(n2913) );
  AOI2BB2XL U9164 ( .B0(n8122), .B1(n7395), .A0N(n9312), .A1N(n8119), .Y(n2789) );
  AOI2BB2XL U9165 ( .B0(n7971), .B1(n7395), .A0N(n9311), .A1N(n7968), .Y(n4639) );
  OA22XL U9166 ( .A0(n7749), .A1(n479), .B0(n8349), .B1(n1107), .Y(n1106) );
  OA22XL U9167 ( .A0(n7741), .A1(n471), .B0(n8349), .B1(n1102), .Y(n1101) );
  OA22XL U9168 ( .A0(n7744), .A1(n857), .B0(n8342), .B1(n1394), .Y(n1393) );
  OA22XL U9169 ( .A0(n7750), .A1(n854), .B0(n8342), .B1(n1390), .Y(n1389) );
  OA22XL U9170 ( .A0(n7745), .A1(n1097), .B0(n8343), .B1(n1625), .Y(n1624) );
  OA22XL U9171 ( .A0(n7745), .A1(n1102), .B0(n8343), .B1(n1628), .Y(n1627) );
  OA22XL U9172 ( .A0(n7746), .A1(n486), .B0(n8346), .B1(n866), .Y(n865) );
  AOI2BB2XL U9173 ( .B0(n7983), .B1(n7393), .A0N(n9326), .A1N(n7979), .Y(n3626) );
  AOI2BB2XL U9174 ( .B0(n8048), .B1(n7393), .A0N(n9324), .A1N(n8044), .Y(n3280) );
  AOI2BB2XL U9175 ( .B0(n8098), .B1(n7393), .A0N(n9322), .A1N(n8095), .Y(n2997) );
  AOI2BB2XL U9176 ( .B0(n8111), .B1(n7393), .A0N(n9321), .A1N(n8107), .Y(n2915) );
  AOI2BB2XL U9177 ( .B0(n8125), .B1(n7393), .A0N(n9320), .A1N(n8121), .Y(n2790) );
  AOI2BB2XL U9178 ( .B0(n7971), .B1(n7393), .A0N(n9319), .A1N(n7967), .Y(n4657) );
  AOI2BB2XL U9179 ( .B0(n7982), .B1(n7391), .A0N(n9334), .A1N(n3572), .Y(n3627) );
  AOI2BB2XL U9180 ( .B0(n8046), .B1(n7391), .A0N(n9332), .A1N(n3226), .Y(n3281) );
  AOI2BB2XL U9181 ( .B0(n8097), .B1(n7391), .A0N(n9330), .A1N(n2943), .Y(n2998) );
  AOI2BB2XL U9182 ( .B0(n8110), .B1(n7391), .A0N(n9329), .A1N(n2808), .Y(n2917) );
  AOI2BB2XL U9183 ( .B0(n8124), .B1(n7391), .A0N(n9328), .A1N(n8119), .Y(n2791) );
  AOI2BB2XL U9184 ( .B0(n7971), .B1(n7391), .A0N(n9327), .A1N(n3654), .Y(n4675) );
  AOI2BB2XL U9185 ( .B0(n7981), .B1(n7389), .A0N(n9342), .A1N(n3572), .Y(n3628) );
  AOI2BB2XL U9186 ( .B0(n8048), .B1(n7389), .A0N(n9340), .A1N(n3226), .Y(n3282) );
  AOI2BB2XL U9187 ( .B0(n8099), .B1(n7389), .A0N(n9338), .A1N(n2943), .Y(n2999) );
  AOI2BB2XL U9188 ( .B0(n8112), .B1(n7389), .A0N(n9337), .A1N(n8106), .Y(n2919) );
  AOI2BB2XL U9189 ( .B0(n8122), .B1(n7389), .A0N(n9336), .A1N(n8121), .Y(n2792) );
  AOI2BB2XL U9190 ( .B0(n7971), .B1(n7389), .A0N(n9335), .A1N(n7966), .Y(n4693) );
  OA22XL U9191 ( .A0(n7749), .A1(n463), .B0(n8348), .B1(n1097), .Y(n1096) );
  OA22XL U9192 ( .A0(n7746), .A1(n851), .B0(n8342), .B1(n1386), .Y(n1385) );
  OA22XL U9193 ( .A0(n7741), .A1(n455), .B0(n8348), .B1(n1092), .Y(n1091) );
  OA22XL U9194 ( .A0(n7750), .A1(n848), .B0(n8342), .B1(n1382), .Y(n1381) );
  OA22XL U9195 ( .A0(n7745), .A1(n1092), .B0(n8343), .B1(n1622), .Y(n1621) );
  OA22XL U9196 ( .A0(n7746), .A1(n462), .B0(n8345), .B1(n857), .Y(n856) );
  AOI2BB2XL U9197 ( .B0(n7981), .B1(n7387), .A0N(n9350), .A1N(n7978), .Y(n3629) );
  AOI2BB2XL U9198 ( .B0(n3225), .B1(n7387), .A0N(n9348), .A1N(n8044), .Y(n3283) );
  AOI2BB2XL U9199 ( .B0(n8097), .B1(n7387), .A0N(n9346), .A1N(n8094), .Y(n3000) );
  AOI2BB2XL U9200 ( .B0(n8109), .B1(n7387), .A0N(n9345), .A1N(n8107), .Y(n2921) );
  AOI2BB2XL U9201 ( .B0(n8122), .B1(n7387), .A0N(n9344), .A1N(n8121), .Y(n2793) );
  AOI2BB2XL U9202 ( .B0(n7971), .B1(n7387), .A0N(n9343), .A1N(n7967), .Y(n4711) );
  AOI2BB2XL U9203 ( .B0(n7984), .B1(n7385), .A0N(n9358), .A1N(n7980), .Y(n3630) );
  AOI2BB2XL U9204 ( .B0(n8045), .B1(n7385), .A0N(n9356), .A1N(n8043), .Y(n3284) );
  AOI2BB2XL U9205 ( .B0(n8096), .B1(n7385), .A0N(n9354), .A1N(n8093), .Y(n3001) );
  AOI2BB2XL U9206 ( .B0(n8109), .B1(n7385), .A0N(n9353), .A1N(n8108), .Y(n2923) );
  AOI2BB2XL U9207 ( .B0(n2735), .B1(n7385), .A0N(n9352), .A1N(n8120), .Y(n2794) );
  AOI2BB2XL U9208 ( .B0(n7971), .B1(n7385), .A0N(n9351), .A1N(n7968), .Y(n4729) );
  AOI2BB2XL U9209 ( .B0(n3571), .B1(n7383), .A0N(n9366), .A1N(n7979), .Y(n3631) );
  AOI2BB2XL U9210 ( .B0(n8047), .B1(n7383), .A0N(n9364), .A1N(n8042), .Y(n3285) );
  AOI2BB2XL U9211 ( .B0(n8096), .B1(n7383), .A0N(n9362), .A1N(n8094), .Y(n3002) );
  AOI2BB2XL U9212 ( .B0(n8110), .B1(n7383), .A0N(n9361), .A1N(n8106), .Y(n2925) );
  AOI2BB2XL U9213 ( .B0(n2735), .B1(n7383), .A0N(n9360), .A1N(n8119), .Y(n2795) );
  AOI2BB2XL U9214 ( .B0(n7971), .B1(n7383), .A0N(n9359), .A1N(n7966), .Y(n4747) );
  OA22XL U9215 ( .A0(n7744), .A1(n470), .B0(n8345), .B1(n860), .Y(n859) );
  OA22XL U9216 ( .A0(n7749), .A1(n447), .B0(n8348), .B1(n1087), .Y(n1086) );
  OA22XL U9217 ( .A0(n7746), .A1(n845), .B0(n8342), .B1(n1378), .Y(n1377) );
  OA22XL U9218 ( .A0(n7741), .A1(n439), .B0(n8348), .B1(n1082), .Y(n1081) );
  OA22XL U9219 ( .A0(n7750), .A1(n842), .B0(n8342), .B1(n1374), .Y(n1373) );
  OA22XL U9220 ( .A0(n7745), .A1(n1087), .B0(n8343), .B1(n1619), .Y(n1618) );
  OA22XL U9221 ( .A0(n7750), .A1(n446), .B0(n8345), .B1(n851), .Y(n850) );
  AOI2BB2XL U9222 ( .B0(n7981), .B1(n7381), .A0N(n9374), .A1N(n7980), .Y(n3632) );
  AOI2BB2XL U9223 ( .B0(n8046), .B1(n7381), .A0N(n9372), .A1N(n8044), .Y(n3286) );
  AOI2BB2XL U9224 ( .B0(n8097), .B1(n7381), .A0N(n9370), .A1N(n2943), .Y(n3003) );
  AOI2BB2XL U9225 ( .B0(n2806), .B1(n7381), .A0N(n9369), .A1N(n8106), .Y(n2927) );
  AOI2BB2XL U9226 ( .B0(n2735), .B1(n7381), .A0N(n9368), .A1N(n8119), .Y(n2796) );
  AOI2BB2XL U9227 ( .B0(n7971), .B1(n7381), .A0N(n9367), .A1N(n3654), .Y(n4765) );
  AOI2BB2XL U9228 ( .B0(n3571), .B1(n7379), .A0N(n9382), .A1N(n3572), .Y(n3633) );
  AOI2BB2XL U9229 ( .B0(n3225), .B1(n7379), .A0N(n9380), .A1N(n8043), .Y(n3287) );
  AOI2BB2XL U9230 ( .B0(n2942), .B1(n7379), .A0N(n9378), .A1N(n8095), .Y(n3004) );
  AOI2BB2XL U9231 ( .B0(n2806), .B1(n7379), .A0N(n9377), .A1N(n8108), .Y(n2929) );
  AOI2BB2XL U9232 ( .B0(n2735), .B1(n7379), .A0N(n9376), .A1N(n8120), .Y(n2797) );
  AOI2BB2XL U9233 ( .B0(n7971), .B1(n7379), .A0N(n9375), .A1N(n7968), .Y(n4783) );
  AOI2BB2XL U9234 ( .B0(n3571), .B1(n7377), .A0N(n9390), .A1N(n7979), .Y(n3634) );
  AOI2BB2XL U9235 ( .B0(n3225), .B1(n7377), .A0N(n9388), .A1N(n3226), .Y(n3288) );
  AOI2BB2XL U9236 ( .B0(n2942), .B1(n7377), .A0N(n9386), .A1N(n8094), .Y(n3005) );
  AOI2BB2XL U9237 ( .B0(n2806), .B1(n7377), .A0N(n9385), .A1N(n2808), .Y(n2931) );
  AOI2BB2XL U9238 ( .B0(n2735), .B1(n7377), .A0N(n9384), .A1N(n8120), .Y(n2798) );
  AOI2BB2XL U9239 ( .B0(n7971), .B1(n7377), .A0N(n9383), .A1N(n7966), .Y(n4801) );
  OA22XL U9240 ( .A0(n7750), .A1(n454), .B0(n8345), .B1(n854), .Y(n853) );
  OA22XL U9241 ( .A0(n7745), .A1(n431), .B0(n8348), .B1(n1077), .Y(n1076) );
  OA22XL U9242 ( .A0(n7744), .A1(n839), .B0(n8342), .B1(n1370), .Y(n1369) );
  OA22XL U9243 ( .A0(n7750), .A1(n836), .B0(n8342), .B1(n1366), .Y(n1365) );
  OA22XL U9244 ( .A0(n7749), .A1(n423), .B0(n8348), .B1(n1072), .Y(n1071) );
  OA22XL U9245 ( .A0(n7741), .A1(n415), .B0(n8348), .B1(n1067), .Y(n1066) );
  OA22XL U9246 ( .A0(n7746), .A1(n833), .B0(n8348), .B1(n1362), .Y(n1361) );
  OA22XL U9247 ( .A0(n7743), .A1(n1077), .B0(n8343), .B1(n1613), .Y(n1612) );
  OA22XL U9248 ( .A0(n7745), .A1(n1072), .B0(n8343), .B1(n1610), .Y(n1609) );
  OA22XL U9249 ( .A0(n7750), .A1(n430), .B0(n8345), .B1(n845), .Y(n844) );
  OA22XL U9250 ( .A0(n7745), .A1(n1067), .B0(n8343), .B1(n1607), .Y(n1606) );
  OA22XL U9251 ( .A0(n7745), .A1(n1062), .B0(n8343), .B1(n1604), .Y(n1603) );
  OA22XL U9252 ( .A0(n7750), .A1(n414), .B0(n8345), .B1(n839), .Y(n838) );
  AOI2BB2XL U9253 ( .B0(n3571), .B1(n7375), .A0N(n9398), .A1N(n7978), .Y(n3635) );
  AOI2BB2XL U9254 ( .B0(n3225), .B1(n7375), .A0N(n9396), .A1N(n8042), .Y(n3289) );
  AOI2BB2XL U9255 ( .B0(n2942), .B1(n7375), .A0N(n9394), .A1N(n8093), .Y(n3006) );
  AOI2BB2XL U9256 ( .B0(n2806), .B1(n7375), .A0N(n9393), .A1N(n8107), .Y(n2933) );
  AOI2BB2XL U9257 ( .B0(n8122), .B1(n7375), .A0N(n9392), .A1N(n8119), .Y(n2799) );
  AOI2BB2XL U9258 ( .B0(n7971), .B1(n7375), .A0N(n9391), .A1N(n7967), .Y(n4819) );
  OA22XL U9259 ( .A0(n7750), .A1(n438), .B0(n8345), .B1(n848), .Y(n847) );
  OA22XL U9260 ( .A0(n7750), .A1(n422), .B0(n8345), .B1(n842), .Y(n841) );
  CLKBUFX2 U9261 ( .A(n8407), .Y(n7227) );
  OA22XL U9262 ( .A0(n7745), .A1(n407), .B0(n8348), .B1(n1062), .Y(n1061) );
  OA22XL U9263 ( .A0(n7745), .A1(n399), .B0(n8348), .B1(n1057), .Y(n1056) );
  OA22XL U9264 ( .A0(n7750), .A1(n830), .B0(n8338), .B1(n1358), .Y(n1357) );
  OA22XL U9265 ( .A0(n7744), .A1(n827), .B0(n8338), .B1(n1354), .Y(n1353) );
  OA22XL U9266 ( .A0(n7754), .A1(n1057), .B0(n8343), .B1(n1601), .Y(n1600) );
  OA22XL U9267 ( .A0(n7754), .A1(n1052), .B0(n8343), .B1(n1598), .Y(n1597) );
  OA22XL U9268 ( .A0(n7741), .A1(n406), .B0(n8345), .B1(n836), .Y(n835) );
  OA22XL U9269 ( .A0(n7758), .A1(n391), .B0(n8348), .B1(n1052), .Y(n1051) );
  OA22XL U9270 ( .A0(n7756), .A1(n383), .B0(n8348), .B1(n1047), .Y(n1046) );
  OA22XL U9271 ( .A0(n7760), .A1(n824), .B0(n8338), .B1(n1350), .Y(n1349) );
  OA22XL U9272 ( .A0(n7760), .A1(n821), .B0(n8342), .B1(n1346), .Y(n1345) );
  OA22XL U9273 ( .A0(n7754), .A1(n1047), .B0(n8343), .B1(n1595), .Y(n1594) );
  OA22XL U9274 ( .A0(n7754), .A1(n1042), .B0(n8343), .B1(n1592), .Y(n1591) );
  OA22XL U9275 ( .A0(n7756), .A1(n390), .B0(n8350), .B1(n830), .Y(n829) );
  OA22XL U9276 ( .A0(n7758), .A1(n375), .B0(n8348), .B1(n1042), .Y(n1041) );
  OA22XL U9277 ( .A0(n7758), .A1(n367), .B0(n8348), .B1(n1037), .Y(n1036) );
  OA22XL U9278 ( .A0(n7760), .A1(n818), .B0(n8339), .B1(n1342), .Y(n1341) );
  OA22XL U9279 ( .A0(n7760), .A1(n815), .B0(n8339), .B1(n1338), .Y(n1337) );
  OA22XL U9280 ( .A0(n7754), .A1(n1037), .B0(n8343), .B1(n1589), .Y(n1588) );
  OA22XL U9281 ( .A0(n7756), .A1(n382), .B0(n8340), .B1(n827), .Y(n826) );
  OA22XL U9282 ( .A0(n7756), .A1(n374), .B0(n8350), .B1(n824), .Y(n823) );
  OA22XL U9283 ( .A0(n7758), .A1(n359), .B0(n8348), .B1(n1032), .Y(n1031) );
  OA22XL U9284 ( .A0(n7758), .A1(n351), .B0(n8348), .B1(n1027), .Y(n1026) );
  OA22XL U9285 ( .A0(n7760), .A1(n812), .B0(n8339), .B1(n1334), .Y(n1333) );
  OA22XL U9286 ( .A0(n7760), .A1(n809), .B0(n8349), .B1(n1330), .Y(n1329) );
  OA22XL U9287 ( .A0(n7754), .A1(n1027), .B0(n8343), .B1(n1583), .Y(n1582) );
  OA22XL U9288 ( .A0(n7756), .A1(n366), .B0(n8340), .B1(n821), .Y(n820) );
  OA22XL U9289 ( .A0(n7754), .A1(n1022), .B0(n8343), .B1(n1580), .Y(n1579) );
  OA22XL U9290 ( .A0(n7756), .A1(n358), .B0(n266), .B1(n818), .Y(n817) );
  OA22XL U9291 ( .A0(n7758), .A1(n343), .B0(n8348), .B1(n1022), .Y(n1021) );
  OA22XL U9292 ( .A0(n7758), .A1(n335), .B0(n8348), .B1(n1017), .Y(n1016) );
  OA22XL U9293 ( .A0(n7760), .A1(n806), .B0(n8337), .B1(n1326), .Y(n1325) );
  OA22XL U9294 ( .A0(n7760), .A1(n803), .B0(n8345), .B1(n1322), .Y(n1321) );
  OA22XL U9295 ( .A0(n7756), .A1(n350), .B0(n266), .B1(n815), .Y(n814) );
  OA22XL U9296 ( .A0(n7754), .A1(n1017), .B0(n8343), .B1(n1577), .Y(n1576) );
  OA22XL U9297 ( .A0(n7754), .A1(n1012), .B0(n8343), .B1(n1574), .Y(n1573) );
  OA22XL U9298 ( .A0(n7756), .A1(n342), .B0(n266), .B1(n812), .Y(n811) );
  OA22XL U9299 ( .A0(n7758), .A1(n327), .B0(n8348), .B1(n1012), .Y(n1011) );
  OA22XL U9300 ( .A0(n7758), .A1(n319), .B0(n8348), .B1(n1007), .Y(n1006) );
  OA22XL U9301 ( .A0(n7760), .A1(n800), .B0(n8345), .B1(n1318), .Y(n1317) );
  OA22XL U9302 ( .A0(n7760), .A1(n797), .B0(n8345), .B1(n1314), .Y(n1313) );
  OA22XL U9303 ( .A0(n7754), .A1(n1007), .B0(n8343), .B1(n1571), .Y(n1570) );
  OA22XL U9304 ( .A0(n7754), .A1(n1002), .B0(n8345), .B1(n1568), .Y(n1567) );
  OA22XL U9305 ( .A0(n7756), .A1(n334), .B0(n266), .B1(n809), .Y(n808) );
  OA22XL U9306 ( .A0(n7756), .A1(n326), .B0(n266), .B1(n806), .Y(n805) );
  OA22XL U9307 ( .A0(n7760), .A1(n794), .B0(n8345), .B1(n1310), .Y(n1309) );
  OA22XL U9308 ( .A0(n7758), .A1(n311), .B0(n8348), .B1(n1002), .Y(n1001) );
  OA22XL U9309 ( .A0(n7754), .A1(n997), .B0(n8345), .B1(n1565), .Y(n1564) );
  OA22XL U9310 ( .A0(n7756), .A1(n318), .B0(n266), .B1(n803), .Y(n802) );
  OA22XL U9311 ( .A0(n7756), .A1(n310), .B0(n8345), .B1(n800), .Y(n799) );
  OA22XL U9312 ( .A0(n7758), .A1(n303), .B0(n8348), .B1(n997), .Y(n996) );
  OA22XL U9313 ( .A0(n7758), .A1(n295), .B0(n8347), .B1(n992), .Y(n991) );
  OA22XL U9314 ( .A0(n7760), .A1(n791), .B0(n8345), .B1(n1306), .Y(n1305) );
  OA22XL U9315 ( .A0(n7754), .A1(n992), .B0(n8345), .B1(n1562), .Y(n1561) );
  OA22XL U9316 ( .A0(n7756), .A1(n294), .B0(n8345), .B1(n794), .Y(n793) );
  OA22XL U9317 ( .A0(n7756), .A1(n302), .B0(n8345), .B1(n797), .Y(n796) );
  OA22XL U9318 ( .A0(n7758), .A1(n287), .B0(n8347), .B1(n987), .Y(n986) );
  OA22XL U9319 ( .A0(n7760), .A1(n788), .B0(n8345), .B1(n1302), .Y(n1301) );
  OA22XL U9320 ( .A0(n7756), .A1(n286), .B0(n8345), .B1(n791), .Y(n790) );
  OA22XL U9321 ( .A0(n7754), .A1(n987), .B0(n8345), .B1(n1559), .Y(n1558) );
  OA22XL U9322 ( .A0(n7758), .A1(n279), .B0(n8347), .B1(n982), .Y(n981) );
  OA22XL U9323 ( .A0(n7754), .A1(n982), .B0(n8345), .B1(n1556), .Y(n1555) );
  OA22XL U9324 ( .A0(n7760), .A1(n784), .B0(n8350), .B1(n1298), .Y(n1297) );
  OA22XL U9325 ( .A0(n7745), .A1(n278), .B0(n8347), .B1(n788), .Y(n787) );
  OA22XL U9326 ( .A0(n7758), .A1(n271), .B0(n8347), .B1(n977), .Y(n976) );
  CLKBUFX3 U9327 ( .A(n2526), .Y(n7502) );
  NAND2X1 U9328 ( .A(n4858), .B(n773), .Y(n4822) );
  NOR2X1 U9329 ( .A(n7002), .B(N1759), .Y(n2524) );
  INVX3 U9330 ( .A(n241), .Y(n8854) );
  NOR2BX1 U9331 ( .AN(n8401), .B(n161), .Y(n160) );
  OA22XL U9332 ( .A0(n7754), .A1(n977), .B0(n8342), .B1(n1553), .Y(n1552) );
  OA22XL U9333 ( .A0(n7745), .A1(n269), .B0(n8341), .B1(n784), .Y(n783) );
  OA22XL U9334 ( .A0(\xArray[1][1] ), .A1(n8187), .B0(\xArray[13][1] ), .B1(
        n8260), .Y(n1740) );
  AOI22XL U9335 ( .A0(n8059), .A1(n7494), .B0(\xArray[8][60] ), .B1(n8055), 
        .Y(n3157) );
  AOI22XL U9336 ( .A0(n8135), .A1(n7494), .B0(\xArray[2][60] ), .B1(n8132), 
        .Y(n2606) );
  AOI22XL U9337 ( .A0(n8059), .A1(n7500), .B0(\xArray[8][63] ), .B1(n8055), 
        .Y(n3152) );
  AOI22XL U9338 ( .A0(n8135), .A1(n7500), .B0(\xArray[2][63] ), .B1(n8132), 
        .Y(n2598) );
  AOI22XL U9339 ( .A0(n8059), .A1(n7496), .B0(\xArray[8][61] ), .B1(n8055), 
        .Y(n3156) );
  AOI22XL U9340 ( .A0(n8135), .A1(n7496), .B0(\xArray[2][61] ), .B1(n8132), 
        .Y(n2604) );
  AOI22XL U9341 ( .A0(n3153), .A1(n7498), .B0(\xArray[8][62] ), .B1(n8055), 
        .Y(n3155) );
  AOI22XL U9342 ( .A0(n8135), .A1(n7498), .B0(\xArray[2][62] ), .B1(n8132), 
        .Y(n2602) );
  NAND2XL U9343 ( .A(n105), .B(n6700), .Y(n779) );
  NAND2XL U9344 ( .A(n6708), .B(n8885), .Y(n775) );
  OA22XL U9345 ( .A0(\xArray[15][1] ), .A1(n8189), .B0(\xArray[11][1] ), .B1(
        n8261), .Y(n2313) );
  OAI221X1 U9346 ( .A0(\xArray[3][1] ), .A1(n8283), .B0(\xArray[7][1] ), .B1(
        n8229), .C0(n2313), .Y(n1546) );
  OA22XL U9347 ( .A0(\xArray[0][1] ), .A1(n8189), .B0(\xArray[12][1] ), .B1(
        n8260), .Y(n2314) );
  OAI221X1 U9348 ( .A0(\xArray[4][1] ), .A1(n8283), .B0(\xArray[8][1] ), .B1(
        n8229), .C0(n2314), .Y(n1544) );
  AOI2BB2XL U9349 ( .B0(n9360), .B1(n8211), .A0N(\xArray[15][4] ), .A1N(n8254), 
        .Y(n1274) );
  OAI221X2 U9350 ( .A0(\xArray[8][2] ), .A1(n8295), .B0(\xArray[12][2] ), .B1(
        n8241), .C0(n1283), .Y(n759) );
  OA22XL U9351 ( .A0(\xArray[4][4] ), .A1(n8198), .B0(\xArray[0][4] ), .B1(
        n8270), .Y(n1273) );
  OA22XL U9352 ( .A0(\xArray[15][2] ), .A1(n8189), .B0(\xArray[11][2] ), .B1(
        n8261), .Y(n2304) );
  OA22XL U9353 ( .A0(\xArray[14][1] ), .A1(n8273), .B0(\xArray[2][1] ), .B1(
        n8187), .Y(n1547) );
  OA22XL U9354 ( .A0(\xArray[1][6] ), .A1(n8187), .B0(\xArray[13][6] ), .B1(
        n8260), .Y(n1725) );
  OA22XL U9355 ( .A0(\xArray[15][0] ), .A1(n8189), .B0(\xArray[11][0] ), .B1(
        n8260), .Y(n2326) );
  AOI22XL U9356 ( .A0(n8059), .A1(n7492), .B0(\xArray[8][59] ), .B1(n8055), 
        .Y(n3158) );
  AOI22XL U9357 ( .A0(n8135), .A1(n7492), .B0(\xArray[2][59] ), .B1(n8132), 
        .Y(n2608) );
  AOI22XL U9358 ( .A0(n8059), .A1(n7490), .B0(\xArray[8][58] ), .B1(n8055), 
        .Y(n3159) );
  AOI22XL U9359 ( .A0(n8135), .A1(n7490), .B0(\xArray[2][58] ), .B1(n8132), 
        .Y(n2610) );
  NAND2XL U9360 ( .A(n103), .B(n8884), .Y(n268) );
  INVXL U9361 ( .A(n104), .Y(n8884) );
  OA22XL U9362 ( .A0(\xArray[14][5] ), .A1(n8272), .B0(\xArray[2][5] ), .B1(
        n8186), .Y(n1531) );
  OAI221X2 U9363 ( .A0(\xArray[9][2] ), .A1(n8290), .B0(\xArray[13][2] ), .B1(
        n8236), .C0(n969), .Y(n758) );
  AND2XL U9364 ( .A(n104), .B(n103), .Y(n6735) );
  AOI2BB2XL U9365 ( .B0(n9358), .B1(n8207), .A0N(\xArray[10][5] ), .A1N(n8258), 
        .Y(n2275) );
  AOI2BB2XL U9366 ( .B0(n9350), .B1(n8208), .A0N(\xArray[10][6] ), .A1N(n8257), 
        .Y(n2266) );
  OA22XL U9367 ( .A0(\xArray[0][7] ), .A1(n8190), .B0(\xArray[12][7] ), .B1(
        n8263), .Y(n2260) );
  OA22XL U9368 ( .A0(\xArray[0][8] ), .A1(n8190), .B0(\xArray[12][8] ), .B1(
        n8263), .Y(n2251) );
  AOI2BB2XL U9369 ( .B0(n9368), .B1(n8210), .A0N(\xArray[15][3] ), .A1N(n8254), 
        .Y(n1279) );
  AOI2BB2XL U9370 ( .B0(n9352), .B1(n8211), .A0N(\xArray[15][5] ), .A1N(n8254), 
        .Y(n1269) );
  OA22XL U9371 ( .A0(\xArray[4][3] ), .A1(n8198), .B0(\xArray[0][3] ), .B1(
        n8270), .Y(n1278) );
  OA22XL U9372 ( .A0(\xArray[4][5] ), .A1(n8198), .B0(\xArray[0][5] ), .B1(
        n8270), .Y(n1268) );
  OA22XL U9373 ( .A0(\xArray[14][7] ), .A1(n8272), .B0(\xArray[2][7] ), .B1(
        n8186), .Y(n1523) );
  OA22XL U9374 ( .A0(\xArray[15][7] ), .A1(n8190), .B0(\xArray[11][7] ), .B1(
        n8263), .Y(n2259) );
  OA22XL U9375 ( .A0(\xArray[15][8] ), .A1(n8190), .B0(\xArray[11][8] ), .B1(
        n8263), .Y(n2250) );
  OA22XL U9376 ( .A0(\xArray[1][7] ), .A1(n8187), .B0(\xArray[13][7] ), .B1(
        n8259), .Y(n1722) );
  AOI22XL U9377 ( .A0(n8059), .A1(n7488), .B0(\xArray[8][57] ), .B1(n8055), 
        .Y(n3160) );
  AOI22XL U9378 ( .A0(n8135), .A1(n7488), .B0(\xArray[2][57] ), .B1(n8132), 
        .Y(n2612) );
  AOI22XL U9379 ( .A0(n8058), .A1(n7486), .B0(\xArray[8][56] ), .B1(n8055), 
        .Y(n3161) );
  AOI22XL U9380 ( .A0(n8135), .A1(n7486), .B0(\xArray[2][56] ), .B1(n8132), 
        .Y(n2614) );
  AOI22XL U9381 ( .A0(n8059), .A1(n7484), .B0(\xArray[8][55] ), .B1(n8055), 
        .Y(n3162) );
  AOI22XL U9382 ( .A0(n8135), .A1(n7484), .B0(\xArray[2][55] ), .B1(n8132), 
        .Y(n2616) );
  OA22XL U9383 ( .A0(\xArray[14][6] ), .A1(n8272), .B0(\xArray[2][6] ), .B1(
        n8186), .Y(n1527) );
  OA22XL U9384 ( .A0(\xArray[5][4] ), .A1(n8196), .B0(\xArray[1][4] ), .B1(
        n8268), .Y(n963) );
  OA22XL U9385 ( .A0(\xArray[5][5] ), .A1(n8196), .B0(\xArray[1][5] ), .B1(
        n8268), .Y(n960) );
  OA22XL U9386 ( .A0(\xArray[5][6] ), .A1(n8196), .B0(\xArray[1][6] ), .B1(
        n8268), .Y(n957) );
  AOI2BB2XL U9387 ( .B0(n9342), .B1(n8208), .A0N(\xArray[10][7] ), .A1N(n8257), 
        .Y(n2257) );
  AOI2BB2XL U9388 ( .B0(n9334), .B1(n8208), .A0N(\xArray[10][8] ), .A1N(n8257), 
        .Y(n2248) );
  AOI2BB2XL U9389 ( .B0(n9344), .B1(n8211), .A0N(\xArray[15][6] ), .A1N(n8254), 
        .Y(n1264) );
  OA22XL U9390 ( .A0(\xArray[4][6] ), .A1(n8198), .B0(\xArray[0][6] ), .B1(
        n8270), .Y(n1263) );
  OA22XL U9391 ( .A0(\xArray[4][7] ), .A1(n8198), .B0(\xArray[0][7] ), .B1(
        n8270), .Y(n1258) );
  OA22XL U9392 ( .A0(\xArray[14][8] ), .A1(n8272), .B0(\xArray[2][8] ), .B1(
        n8186), .Y(n1519) );
  OA22XL U9393 ( .A0(\xArray[14][9] ), .A1(n8273), .B0(\xArray[2][9] ), .B1(
        n8186), .Y(n1515) );
  OA22XL U9394 ( .A0(\xArray[1][8] ), .A1(n8187), .B0(\xArray[13][8] ), .B1(
        n8260), .Y(n1719) );
  OA22XL U9395 ( .A0(\xArray[1][9] ), .A1(n8187), .B0(\xArray[13][9] ), .B1(
        n8259), .Y(n1716) );
  AOI22XL U9396 ( .A0(n8060), .A1(n7482), .B0(\xArray[8][54] ), .B1(n8055), 
        .Y(n3163) );
  AOI22XL U9397 ( .A0(n8135), .A1(n7482), .B0(\xArray[2][54] ), .B1(n8132), 
        .Y(n2618) );
  AOI22XL U9398 ( .A0(n3153), .A1(n7480), .B0(\xArray[8][53] ), .B1(n8055), 
        .Y(n3164) );
  AOI22XL U9399 ( .A0(n8135), .A1(n7480), .B0(\xArray[2][53] ), .B1(n8132), 
        .Y(n2620) );
  AOI22XL U9400 ( .A0(n8059), .A1(n7478), .B0(\xArray[8][52] ), .B1(n8055), 
        .Y(n3165) );
  AOI22XL U9401 ( .A0(n8135), .A1(n7478), .B0(\xArray[2][52] ), .B1(n8132), 
        .Y(n2622) );
  AOI2BB2XL U9402 ( .B0(n9336), .B1(n8211), .A0N(\xArray[15][7] ), .A1N(n8254), 
        .Y(n1259) );
  INVXL U9403 ( .A(\xArray[3][4] ), .Y(n9360) );
  OA22XL U9404 ( .A0(n8321), .A1(n1550), .B0(n7728), .B1(n1742), .Y(n2315) );
  OA22XL U9405 ( .A0(\xArray[5][7] ), .A1(n8196), .B0(\xArray[1][7] ), .B1(
        n8268), .Y(n954) );
  OA22XL U9406 ( .A0(\xArray[5][8] ), .A1(n8196), .B0(\xArray[1][8] ), .B1(
        n8268), .Y(n951) );
  AOI2BB2XL U9407 ( .B0(n9326), .B1(n8208), .A0N(\xArray[10][9] ), .A1N(n8257), 
        .Y(n2239) );
  AOI2BB2XL U9408 ( .B0(n9318), .B1(n8208), .A0N(\xArray[10][10] ), .A1N(n8258), .Y(n2230) );
  OA22XL U9409 ( .A0(\xArray[4][9] ), .A1(n8198), .B0(\xArray[0][9] ), .B1(
        n8270), .Y(n1248) );
  OA22XL U9410 ( .A0(\xArray[14][11] ), .A1(n8272), .B0(\xArray[2][11] ), .B1(
        n8186), .Y(n1507) );
  OA22XL U9411 ( .A0(\xArray[1][10] ), .A1(n8187), .B0(\xArray[13][10] ), .B1(
        n8259), .Y(n1713) );
  OA22XL U9412 ( .A0(\xArray[1][11] ), .A1(n8187), .B0(\xArray[13][11] ), .B1(
        n8260), .Y(n1710) );
  AOI22XL U9413 ( .A0(n8059), .A1(n7476), .B0(\xArray[8][51] ), .B1(n8055), 
        .Y(n3166) );
  AOI22XL U9414 ( .A0(n8136), .A1(n7476), .B0(\xArray[2][51] ), .B1(n8133), 
        .Y(n2624) );
  AOI22XL U9415 ( .A0(n8059), .A1(n7474), .B0(\xArray[8][50] ), .B1(n8057), 
        .Y(n3167) );
  AOI22XL U9416 ( .A0(n8136), .A1(n7474), .B0(\xArray[2][50] ), .B1(n8133), 
        .Y(n2626) );
  AOI22XL U9417 ( .A0(n8059), .A1(n7472), .B0(\xArray[8][49] ), .B1(n8055), 
        .Y(n3168) );
  AOI22XL U9418 ( .A0(n8136), .A1(n7472), .B0(\xArray[2][49] ), .B1(n8133), 
        .Y(n2628) );
  OA22XL U9419 ( .A0(n8323), .A1(n1538), .B0(n7728), .B1(n1733), .Y(n2288) );
  INVXL U9420 ( .A(\xArray[14][7] ), .Y(n9342) );
  AOI2BB2XL U9421 ( .B0(n9328), .B1(n8211), .A0N(\xArray[15][8] ), .A1N(n8254), 
        .Y(n1254) );
  AOI2BB2XL U9422 ( .B0(n9320), .B1(n8211), .A0N(\xArray[15][9] ), .A1N(n8254), 
        .Y(n1249) );
  INVXL U9423 ( .A(\xArray[3][5] ), .Y(n9352) );
  INVXL U9424 ( .A(\xArray[3][6] ), .Y(n9344) );
  OA22XL U9425 ( .A0(\xArray[5][9] ), .A1(n8196), .B0(\xArray[1][9] ), .B1(
        n8268), .Y(n948) );
  OA22XL U9426 ( .A0(\xArray[5][10] ), .A1(n8196), .B0(\xArray[1][10] ), .B1(
        n8269), .Y(n945) );
  AOI2BB2XL U9427 ( .B0(n9310), .B1(n8208), .A0N(\xArray[10][11] ), .A1N(n8258), .Y(n2221) );
  OA22XL U9428 ( .A0(\xArray[0][12] ), .A1(n8190), .B0(\xArray[12][12] ), .B1(
        n8264), .Y(n2215) );
  OA22XL U9429 ( .A0(\xArray[0][13] ), .A1(n8190), .B0(\xArray[12][13] ), .B1(
        n8264), .Y(n2206) );
  OA22XL U9430 ( .A0(\xArray[1][12] ), .A1(n8187), .B0(\xArray[13][12] ), .B1(
        n8259), .Y(n1707) );
  OA22XL U9431 ( .A0(\xArray[4][10] ), .A1(n8198), .B0(\xArray[0][10] ), .B1(
        n8270), .Y(n1243) );
  OA22XL U9432 ( .A0(\xArray[4][11] ), .A1(n8198), .B0(\xArray[0][11] ), .B1(
        n8270), .Y(n1238) );
  OA22XL U9433 ( .A0(\xArray[14][12] ), .A1(n8272), .B0(\xArray[2][12] ), .B1(
        n8186), .Y(n1503) );
  OA22XL U9434 ( .A0(\xArray[14][13] ), .A1(n8272), .B0(\xArray[2][13] ), .B1(
        n8186), .Y(n1499) );
  OA22XL U9435 ( .A0(\xArray[1][13] ), .A1(n8187), .B0(\xArray[13][13] ), .B1(
        n8259), .Y(n1704) );
  AOI22XL U9436 ( .A0(n8059), .A1(n7470), .B0(\xArray[8][48] ), .B1(n8056), 
        .Y(n3169) );
  AOI22XL U9437 ( .A0(n8136), .A1(n7470), .B0(\xArray[2][48] ), .B1(n8133), 
        .Y(n2630) );
  AOI22XL U9438 ( .A0(n8059), .A1(n7468), .B0(\xArray[8][47] ), .B1(n8057), 
        .Y(n3170) );
  AOI22XL U9439 ( .A0(n8136), .A1(n7468), .B0(\xArray[2][47] ), .B1(n8133), 
        .Y(n2632) );
  AOI22XL U9440 ( .A0(n8059), .A1(n7466), .B0(\xArray[8][46] ), .B1(n8055), 
        .Y(n3171) );
  AOI22XL U9441 ( .A0(n8136), .A1(n7466), .B0(\xArray[2][46] ), .B1(n8133), 
        .Y(n2634) );
  OA22XL U9442 ( .A0(n8323), .A1(n1534), .B0(n7728), .B1(n1730), .Y(n2279) );
  OA22XL U9443 ( .A0(n8323), .A1(n1530), .B0(n7728), .B1(n1727), .Y(n2270) );
  INVXL U9444 ( .A(\xArray[14][8] ), .Y(n9334) );
  INVXL U9445 ( .A(\xArray[14][9] ), .Y(n9326) );
  AOI2BB2XL U9446 ( .B0(n9312), .B1(n8211), .A0N(\xArray[15][10] ), .A1N(n8254), .Y(n1244) );
  INVXL U9447 ( .A(\xArray[3][7] ), .Y(n9336) );
  INVXL U9448 ( .A(\xArray[3][8] ), .Y(n9328) );
  OA22XL U9449 ( .A0(\xArray[15][12] ), .A1(n8190), .B0(\xArray[11][12] ), 
        .B1(n8264), .Y(n2214) );
  OA22XL U9450 ( .A0(\xArray[15][13] ), .A1(n8190), .B0(\xArray[11][13] ), 
        .B1(n8264), .Y(n2205) );
  AOI2BB2XL U9451 ( .B0(n9302), .B1(n8208), .A0N(\xArray[10][12] ), .A1N(n8258), .Y(n2212) );
  OA22XL U9452 ( .A0(\xArray[5][11] ), .A1(n8196), .B0(\xArray[1][11] ), .B1(
        n8269), .Y(n942) );
  OA22XL U9453 ( .A0(\xArray[5][12] ), .A1(n8196), .B0(\xArray[1][12] ), .B1(
        n8269), .Y(n939) );
  AOI2BB2XL U9454 ( .B0(n9294), .B1(n8209), .A0N(\xArray[10][13] ), .A1N(n8258), .Y(n2203) );
  AOI2BB2XL U9455 ( .B0(n9286), .B1(n8209), .A0N(\xArray[10][14] ), .A1N(n8258), .Y(n2194) );
  OA22XL U9456 ( .A0(\xArray[0][15] ), .A1(n8190), .B0(\xArray[12][15] ), .B1(
        n8265), .Y(n2188) );
  OA22XL U9457 ( .A0(\xArray[0][14] ), .A1(n8190), .B0(\xArray[12][14] ), .B1(
        n8264), .Y(n2197) );
  OA22XL U9458 ( .A0(\xArray[4][12] ), .A1(n8198), .B0(\xArray[0][12] ), .B1(
        n8270), .Y(n1233) );
  OA22XL U9459 ( .A0(\xArray[4][13] ), .A1(n8198), .B0(\xArray[0][13] ), .B1(
        n8270), .Y(n1228) );
  OA22XL U9460 ( .A0(\xArray[14][14] ), .A1(n8271), .B0(\xArray[2][14] ), .B1(
        n8186), .Y(n1495) );
  OA22XL U9461 ( .A0(\xArray[14][15] ), .A1(n8272), .B0(\xArray[2][15] ), .B1(
        n8186), .Y(n1491) );
  AOI22XL U9462 ( .A0(n8059), .A1(n7464), .B0(\xArray[8][45] ), .B1(n8056), 
        .Y(n3172) );
  AOI22XL U9463 ( .A0(n8136), .A1(n7464), .B0(\xArray[2][45] ), .B1(n8133), 
        .Y(n2636) );
  AOI22XL U9464 ( .A0(n8059), .A1(n7462), .B0(\xArray[8][44] ), .B1(n8057), 
        .Y(n3173) );
  AOI22XL U9465 ( .A0(n8136), .A1(n7462), .B0(\xArray[2][44] ), .B1(n8133), 
        .Y(n2638) );
  OA22XL U9466 ( .A0(n8323), .A1(n1526), .B0(n7728), .B1(n1724), .Y(n2261) );
  OA22XL U9467 ( .A0(n8323), .A1(n1522), .B0(n7728), .B1(n1721), .Y(n2252) );
  INVXL U9468 ( .A(\xArray[14][10] ), .Y(n9318) );
  INVXL U9469 ( .A(\xArray[14][11] ), .Y(n9310) );
  INVXL U9470 ( .A(\xArray[5][1] ), .Y(n9386) );
  INVXL U9471 ( .A(\xArray[5][0] ), .Y(n9394) );
  INVXL U9472 ( .A(\xArray[5][2] ), .Y(n9378) );
  INVXL U9473 ( .A(\xArray[3][9] ), .Y(n9320) );
  INVXL U9474 ( .A(\xArray[3][10] ), .Y(n9312) );
  INVXL U9475 ( .A(\xArray[9][1] ), .Y(n9388) );
  INVXL U9476 ( .A(\xArray[9][0] ), .Y(n9396) );
  INVXL U9477 ( .A(\xArray[9][2] ), .Y(n9380) );
  INVXL U9478 ( .A(\xArray[6][0] ), .Y(n9395) );
  INVXL U9479 ( .A(\xArray[6][1] ), .Y(n9387) );
  INVXL U9480 ( .A(\xArray[10][0] ), .Y(n9397) );
  INVXL U9481 ( .A(\xArray[10][1] ), .Y(n9389) );
  OA22XL U9482 ( .A0(\xArray[15][15] ), .A1(n8190), .B0(\xArray[11][15] ), 
        .B1(n8265), .Y(n2187) );
  OA22XL U9483 ( .A0(\xArray[15][14] ), .A1(n8190), .B0(\xArray[11][14] ), 
        .B1(n8264), .Y(n2196) );
  OA22XL U9484 ( .A0(\xArray[5][13] ), .A1(n8196), .B0(\xArray[1][13] ), .B1(
        n8269), .Y(n936) );
  OA22XL U9485 ( .A0(\xArray[5][14] ), .A1(n8196), .B0(\xArray[1][14] ), .B1(
        n8269), .Y(n933) );
  AOI2BB2XL U9486 ( .B0(n9278), .B1(n8209), .A0N(\xArray[10][15] ), .A1N(n8258), .Y(n2185) );
  AOI2BB2XL U9487 ( .B0(n9270), .B1(n8209), .A0N(\xArray[10][16] ), .A1N(n8258), .Y(n2176) );
  OA22XL U9488 ( .A0(\xArray[0][16] ), .A1(n8190), .B0(\xArray[12][16] ), .B1(
        n8265), .Y(n2179) );
  OA22XL U9489 ( .A0(\xArray[14][17] ), .A1(n8272), .B0(\xArray[2][17] ), .B1(
        n8186), .Y(n1483) );
  OA22XL U9490 ( .A0(\xArray[4][14] ), .A1(n8198), .B0(\xArray[0][14] ), .B1(
        n8270), .Y(n1223) );
  OA22XL U9491 ( .A0(\xArray[4][15] ), .A1(n8198), .B0(\xArray[0][15] ), .B1(
        n8268), .Y(n1218) );
  OA22XL U9492 ( .A0(\xArray[14][16] ), .A1(n8271), .B0(\xArray[2][16] ), .B1(
        n8186), .Y(n1487) );
  OA22XL U9493 ( .A0(\xArray[1][17] ), .A1(n8188), .B0(\xArray[13][17] ), .B1(
        n8260), .Y(n1692) );
  AOI22XL U9494 ( .A0(n8059), .A1(n7461), .B0(\xArray[8][43] ), .B1(n8055), 
        .Y(n3174) );
  AOI22XL U9495 ( .A0(n8136), .A1(n7461), .B0(\xArray[2][43] ), .B1(n8133), 
        .Y(n2640) );
  AOI22XL U9496 ( .A0(n8059), .A1(n7459), .B0(\xArray[8][42] ), .B1(n3154), 
        .Y(n3175) );
  AOI22XL U9497 ( .A0(n8136), .A1(n7459), .B0(\xArray[2][42] ), .B1(n8133), 
        .Y(n2642) );
  AOI22XL U9498 ( .A0(n8059), .A1(n7457), .B0(\xArray[8][41] ), .B1(n8056), 
        .Y(n3176) );
  AOI22XL U9499 ( .A0(n8136), .A1(n7457), .B0(\xArray[2][41] ), .B1(n8133), 
        .Y(n2644) );
  OA22XL U9500 ( .A0(n8322), .A1(n1518), .B0(n7728), .B1(n1718), .Y(n2243) );
  OA22XL U9501 ( .A0(n8322), .A1(n1514), .B0(n7728), .B1(n1715), .Y(n2234) );
  INVXL U9502 ( .A(\xArray[14][12] ), .Y(n9302) );
  INVXL U9503 ( .A(\xArray[14][13] ), .Y(n9294) );
  INVXL U9504 ( .A(\xArray[5][3] ), .Y(n9370) );
  INVXL U9505 ( .A(\xArray[3][11] ), .Y(n9304) );
  INVXL U9506 ( .A(\xArray[3][12] ), .Y(n9296) );
  INVXL U9507 ( .A(\xArray[9][3] ), .Y(n9372) );
  INVXL U9508 ( .A(\xArray[6][2] ), .Y(n9379) );
  INVXL U9509 ( .A(\xArray[6][3] ), .Y(n9371) );
  INVXL U9510 ( .A(\xArray[10][2] ), .Y(n9381) );
  INVXL U9511 ( .A(\xArray[10][3] ), .Y(n9373) );
  OA22XL U9512 ( .A0(\xArray[5][15] ), .A1(n8196), .B0(\xArray[1][15] ), .B1(
        n8269), .Y(n930) );
  AOI2BB2XL U9513 ( .B0(n9262), .B1(n8209), .A0N(\xArray[10][17] ), .A1N(n8258), .Y(n2167) );
  AOI2BB2XL U9514 ( .B0(n9254), .B1(n8209), .A0N(\xArray[10][18] ), .A1N(n8258), .Y(n2158) );
  OA22XL U9515 ( .A0(\xArray[4][16] ), .A1(n8198), .B0(\xArray[0][16] ), .B1(
        n8267), .Y(n1213) );
  OA22XL U9516 ( .A0(\xArray[14][18] ), .A1(n8271), .B0(\xArray[2][18] ), .B1(
        n8186), .Y(n1479) );
  OA22XL U9517 ( .A0(\xArray[14][19] ), .A1(n8272), .B0(\xArray[2][19] ), .B1(
        n8186), .Y(n1475) );
  OA22XL U9518 ( .A0(\xArray[1][19] ), .A1(n8188), .B0(\xArray[13][19] ), .B1(
        n8261), .Y(n1686) );
  AOI22XL U9519 ( .A0(n8059), .A1(n7455), .B0(\xArray[8][40] ), .B1(n8055), 
        .Y(n3177) );
  AOI22XL U9520 ( .A0(n8136), .A1(n7455), .B0(\xArray[2][40] ), .B1(n8133), 
        .Y(n2646) );
  AOI22XL U9521 ( .A0(n8058), .A1(n7453), .B0(\xArray[8][39] ), .B1(n8056), 
        .Y(n3178) );
  AOI22XL U9522 ( .A0(n8135), .A1(n7453), .B0(\xArray[2][39] ), .B1(n2601), 
        .Y(n2648) );
  AOI22XL U9523 ( .A0(n8058), .A1(n7451), .B0(\xArray[8][38] ), .B1(n8056), 
        .Y(n3179) );
  AOI22XL U9524 ( .A0(n8136), .A1(n7451), .B0(\xArray[2][38] ), .B1(n8134), 
        .Y(n2650) );
  OA22XL U9525 ( .A0(n8322), .A1(n1510), .B0(n7728), .B1(n1712), .Y(n2225) );
  INVXL U9526 ( .A(\xArray[14][14] ), .Y(n9286) );
  INVXL U9527 ( .A(\xArray[14][15] ), .Y(n9278) );
  INVXL U9528 ( .A(\xArray[5][4] ), .Y(n9362) );
  INVXL U9529 ( .A(\xArray[5][5] ), .Y(n9354) );
  INVXL U9530 ( .A(\xArray[3][13] ), .Y(n9288) );
  INVXL U9531 ( .A(\xArray[3][14] ), .Y(n9280) );
  INVXL U9532 ( .A(\xArray[9][4] ), .Y(n9364) );
  INVXL U9533 ( .A(\xArray[9][5] ), .Y(n9356) );
  INVXL U9534 ( .A(\xArray[6][4] ), .Y(n9363) );
  INVXL U9535 ( .A(\xArray[10][4] ), .Y(n9365) );
  INVXL U9536 ( .A(\xArray[10][5] ), .Y(n9357) );
  AOI2BB2XL U9537 ( .B0(n9246), .B1(n8209), .A0N(\xArray[10][19] ), .A1N(n8258), .Y(n2149) );
  AOI2BB2XL U9538 ( .B0(n9238), .B1(n8210), .A0N(\xArray[10][20] ), .A1N(n8258), .Y(n2140) );
  AOI2BB2XL U9539 ( .B0(n9248), .B1(n8208), .A0N(\xArray[15][18] ), .A1N(n8255), .Y(n1204) );
  AOI2BB2XL U9540 ( .B0(n9240), .B1(n8207), .A0N(\xArray[15][19] ), .A1N(n8255), .Y(n1199) );
  OA22XL U9541 ( .A0(\xArray[4][18] ), .A1(n8197), .B0(\xArray[0][18] ), .B1(
        n8267), .Y(n1203) );
  OA22XL U9542 ( .A0(\xArray[4][19] ), .A1(n8197), .B0(\xArray[0][19] ), .B1(
        n8267), .Y(n1198) );
  OA22XL U9543 ( .A0(\xArray[14][21] ), .A1(n8272), .B0(\xArray[2][21] ), .B1(
        n8186), .Y(n1467) );
  OA22XL U9544 ( .A0(\xArray[14][20] ), .A1(n8271), .B0(\xArray[2][20] ), .B1(
        n8186), .Y(n1471) );
  OA22XL U9545 ( .A0(\xArray[1][21] ), .A1(n8188), .B0(\xArray[13][21] ), .B1(
        n8260), .Y(n1680) );
  OA22XL U9546 ( .A0(\xArray[1][20] ), .A1(n8188), .B0(\xArray[13][20] ), .B1(
        n8260), .Y(n1683) );
  AOI22XL U9547 ( .A0(n8058), .A1(n7449), .B0(\xArray[8][37] ), .B1(n8056), 
        .Y(n3180) );
  AOI22XL U9548 ( .A0(n8135), .A1(n7449), .B0(\xArray[2][37] ), .B1(n8132), 
        .Y(n2652) );
  AOI22XL U9549 ( .A0(n8058), .A1(n7447), .B0(\xArray[8][36] ), .B1(n8056), 
        .Y(n3181) );
  AOI22XL U9550 ( .A0(n8136), .A1(n7447), .B0(\xArray[2][36] ), .B1(n8133), 
        .Y(n2654) );
  AOI22XL U9551 ( .A0(n8058), .A1(n7445), .B0(\xArray[8][35] ), .B1(n8056), 
        .Y(n3182) );
  AOI22XL U9552 ( .A0(n8135), .A1(n7445), .B0(\xArray[2][35] ), .B1(n8134), 
        .Y(n2656) );
  INVXL U9553 ( .A(\xArray[14][16] ), .Y(n9270) );
  INVXL U9554 ( .A(\xArray[14][17] ), .Y(n9262) );
  INVXL U9555 ( .A(\xArray[5][6] ), .Y(n9346) );
  INVXL U9556 ( .A(\xArray[5][7] ), .Y(n9338) );
  INVXL U9557 ( .A(\xArray[3][15] ), .Y(n9272) );
  INVXL U9558 ( .A(\xArray[9][6] ), .Y(n9348) );
  INVXL U9559 ( .A(\xArray[9][7] ), .Y(n9340) );
  INVXL U9560 ( .A(\xArray[6][5] ), .Y(n9355) );
  INVXL U9561 ( .A(\xArray[6][6] ), .Y(n9347) );
  INVXL U9562 ( .A(\xArray[10][6] ), .Y(n9349) );
  OA22XL U9563 ( .A0(\xArray[5][20] ), .A1(n8195), .B0(\xArray[1][20] ), .B1(
        n8269), .Y(n915) );
  AOI2BB2XL U9564 ( .B0(n9230), .B1(n8210), .A0N(\xArray[10][21] ), .A1N(n8258), .Y(n2131) );
  AOI2BB2XL U9565 ( .B0(n9232), .B1(n8208), .A0N(\xArray[15][20] ), .A1N(n8255), .Y(n1194) );
  AOI2BB2XL U9566 ( .B0(n9224), .B1(n8208), .A0N(\xArray[15][21] ), .A1N(n8255), .Y(n1189) );
  OA22XL U9567 ( .A0(\xArray[1][22] ), .A1(n8188), .B0(\xArray[13][22] ), .B1(
        n8261), .Y(n1677) );
  OA22XL U9568 ( .A0(\xArray[4][20] ), .A1(n8197), .B0(\xArray[0][20] ), .B1(
        n8267), .Y(n1193) );
  OA22XL U9569 ( .A0(\xArray[4][21] ), .A1(n8197), .B0(\xArray[0][21] ), .B1(
        n8267), .Y(n1188) );
  OA22XL U9570 ( .A0(\xArray[14][22] ), .A1(n8271), .B0(\xArray[2][22] ), .B1(
        n8186), .Y(n1463) );
  AOI22XL U9571 ( .A0(n8058), .A1(n7443), .B0(\xArray[8][34] ), .B1(n8056), 
        .Y(n3183) );
  AOI22XL U9572 ( .A0(n8136), .A1(n7443), .B0(\xArray[2][34] ), .B1(n8132), 
        .Y(n2658) );
  AOI22XL U9573 ( .A0(n8058), .A1(n7441), .B0(\xArray[8][33] ), .B1(n8056), 
        .Y(n3184) );
  AOI22XL U9574 ( .A0(n8137), .A1(n7441), .B0(\xArray[2][33] ), .B1(n8133), 
        .Y(n2660) );
  AOI22XL U9575 ( .A0(n8060), .A1(n7439), .B0(\xArray[8][32] ), .B1(n8056), 
        .Y(n3185) );
  AOI22XL U9576 ( .A0(n8135), .A1(n7439), .B0(\xArray[2][32] ), .B1(n8133), 
        .Y(n2662) );
  MX4XL U9577 ( .A(\bArray[4][17] ), .B(\bArray[5][17] ), .C(\bArray[6][17] ), 
        .D(\bArray[7][17] ), .S0(n7205), .S1(n7217), .Y(n7014) );
  MX4XL U9578 ( .A(\bArray[12][17] ), .B(\bArray[13][17] ), .C(
        \bArray[14][17] ), .D(\bArray[15][17] ), .S0(n7205), .S1(n7217), .Y(
        n7012) );
  MX4XL U9579 ( .A(\bArray[8][17] ), .B(\bArray[9][17] ), .C(\bArray[10][17] ), 
        .D(\bArray[11][17] ), .S0(n7205), .S1(n7217), .Y(n7013) );
  MX4XL U9580 ( .A(\bArray[12][18] ), .B(\bArray[13][18] ), .C(
        \bArray[14][18] ), .D(\bArray[15][18] ), .S0(n7205), .S1(n7217), .Y(
        n7016) );
  MX4XL U9581 ( .A(\bArray[8][18] ), .B(\bArray[9][18] ), .C(\bArray[10][18] ), 
        .D(\bArray[11][18] ), .S0(n7205), .S1(n7217), .Y(n7017) );
  MX4XL U9582 ( .A(\bArray[4][19] ), .B(\bArray[5][19] ), .C(\bArray[6][19] ), 
        .D(\bArray[7][19] ), .S0(n7206), .S1(n7218), .Y(n7022) );
  MX4XL U9583 ( .A(\bArray[12][19] ), .B(\bArray[13][19] ), .C(
        \bArray[14][19] ), .D(\bArray[15][19] ), .S0(n7206), .S1(n7218), .Y(
        n7020) );
  MX4XL U9584 ( .A(\bArray[8][19] ), .B(\bArray[9][19] ), .C(\bArray[10][19] ), 
        .D(\bArray[11][19] ), .S0(n7206), .S1(n7218), .Y(n7021) );
  INVXL U9585 ( .A(\xArray[14][18] ), .Y(n9254) );
  INVXL U9586 ( .A(\xArray[5][8] ), .Y(n9330) );
  INVXL U9587 ( .A(\xArray[5][9] ), .Y(n9322) );
  INVXL U9588 ( .A(\xArray[3][16] ), .Y(n9264) );
  INVXL U9589 ( .A(\xArray[3][17] ), .Y(n9256) );
  INVXL U9590 ( .A(\xArray[9][8] ), .Y(n9332) );
  INVXL U9591 ( .A(\xArray[9][9] ), .Y(n9324) );
  INVXL U9592 ( .A(\xArray[6][7] ), .Y(n9339) );
  INVXL U9593 ( .A(\xArray[6][8] ), .Y(n9331) );
  INVXL U9594 ( .A(\xArray[10][7] ), .Y(n9341) );
  INVXL U9595 ( .A(\xArray[10][8] ), .Y(n9333) );
  MX4XL U9596 ( .A(\bArray[0][17] ), .B(\bArray[1][17] ), .C(\bArray[2][17] ), 
        .D(\bArray[3][17] ), .S0(n7205), .S1(n7217), .Y(n7015) );
  AOI2BB2XL U9597 ( .B0(n9222), .B1(n8210), .A0N(\xArray[10][22] ), .A1N(n8259), .Y(n2122) );
  OA22XL U9598 ( .A0(\xArray[5][21] ), .A1(n8195), .B0(\xArray[1][21] ), .B1(
        n8269), .Y(n912) );
  OA22XL U9599 ( .A0(\xArray[5][22] ), .A1(n8195), .B0(\xArray[1][22] ), .B1(
        n8269), .Y(n909) );
  AOI2BB2XL U9600 ( .B0(n9214), .B1(n8210), .A0N(\xArray[10][23] ), .A1N(n8259), .Y(n2113) );
  OA22XL U9601 ( .A0(\xArray[0][25] ), .A1(n8191), .B0(\xArray[12][25] ), .B1(
        n8267), .Y(n2098) );
  OA22XL U9602 ( .A0(\xArray[0][24] ), .A1(n8191), .B0(\xArray[12][24] ), .B1(
        n8266), .Y(n2107) );
  AOI2BB2XL U9603 ( .B0(n9216), .B1(n8207), .A0N(\xArray[15][22] ), .A1N(n8255), .Y(n1184) );
  OA22XL U9604 ( .A0(\xArray[4][23] ), .A1(n8197), .B0(\xArray[0][23] ), .B1(
        n8267), .Y(n1178) );
  OA22XL U9605 ( .A0(\xArray[4][22] ), .A1(n8197), .B0(\xArray[0][22] ), .B1(
        n8267), .Y(n1183) );
  OA22XL U9606 ( .A0(\xArray[14][24] ), .A1(n8271), .B0(\xArray[2][24] ), .B1(
        n8186), .Y(n1455) );
  OA22XL U9607 ( .A0(\xArray[14][23] ), .A1(n8271), .B0(\xArray[2][23] ), .B1(
        n8186), .Y(n1459) );
  OA22XL U9608 ( .A0(\xArray[15][25] ), .A1(n8191), .B0(\xArray[11][25] ), 
        .B1(n8263), .Y(n2097) );
  OA22XL U9609 ( .A0(\xArray[15][24] ), .A1(n8191), .B0(\xArray[11][24] ), 
        .B1(n8266), .Y(n2106) );
  OA22XL U9610 ( .A0(\xArray[1][24] ), .A1(n8188), .B0(\xArray[13][24] ), .B1(
        n8261), .Y(n1671) );
  AOI22XL U9611 ( .A0(n8060), .A1(n7437), .B0(\xArray[8][31] ), .B1(n8056), 
        .Y(n3186) );
  AOI22XL U9612 ( .A0(n8135), .A1(n7437), .B0(\xArray[2][31] ), .B1(n8133), 
        .Y(n2664) );
  AOI22XL U9613 ( .A0(n8058), .A1(n7435), .B0(\xArray[8][30] ), .B1(n8056), 
        .Y(n3187) );
  AOI22XL U9614 ( .A0(n2599), .A1(n7435), .B0(\xArray[2][30] ), .B1(n8134), 
        .Y(n2666) );
  AOI22XL U9615 ( .A0(n8058), .A1(n7433), .B0(\xArray[8][29] ), .B1(n8056), 
        .Y(n3188) );
  AOI22XL U9616 ( .A0(n2599), .A1(n7433), .B0(\xArray[2][29] ), .B1(n8132), 
        .Y(n2668) );
  OA22XL U9617 ( .A0(n8322), .A1(n1482), .B0(n7729), .B1(n1691), .Y(n2162) );
  OA22XL U9618 ( .A0(n8322), .A1(n1486), .B0(n7729), .B1(n1694), .Y(n2171) );
  MX4XL U9619 ( .A(\bArray[4][20] ), .B(\bArray[5][20] ), .C(\bArray[6][20] ), 
        .D(\bArray[7][20] ), .S0(n7206), .S1(n7218), .Y(n7026) );
  MX4XL U9620 ( .A(\bArray[12][20] ), .B(\bArray[13][20] ), .C(
        \bArray[14][20] ), .D(\bArray[15][20] ), .S0(n7206), .S1(n7218), .Y(
        n7024) );
  MX4XL U9621 ( .A(\bArray[8][20] ), .B(\bArray[9][20] ), .C(\bArray[10][20] ), 
        .D(\bArray[11][20] ), .S0(n7206), .S1(n7218), .Y(n7025) );
  INVXL U9622 ( .A(\xArray[14][19] ), .Y(n9246) );
  INVXL U9623 ( .A(\xArray[14][20] ), .Y(n9238) );
  INVXL U9624 ( .A(\xArray[5][10] ), .Y(n9314) );
  INVXL U9625 ( .A(\xArray[5][11] ), .Y(n9306) );
  INVXL U9626 ( .A(\xArray[3][18] ), .Y(n9248) );
  INVXL U9627 ( .A(\xArray[3][19] ), .Y(n9240) );
  INVXL U9628 ( .A(\xArray[9][10] ), .Y(n9316) );
  INVXL U9629 ( .A(\xArray[9][11] ), .Y(n9308) );
  INVXL U9630 ( .A(\xArray[6][9] ), .Y(n9323) );
  INVXL U9631 ( .A(\xArray[6][10] ), .Y(n9315) );
  INVXL U9632 ( .A(\xArray[10][9] ), .Y(n9325) );
  INVXL U9633 ( .A(\xArray[10][10] ), .Y(n9317) );
  MX4XL U9634 ( .A(\bArray[0][19] ), .B(\bArray[1][19] ), .C(\bArray[2][19] ), 
        .D(\bArray[3][19] ), .S0(n7206), .S1(n7218), .Y(n7023) );
  MX4XL U9635 ( .A(\bArray[0][20] ), .B(\bArray[1][20] ), .C(\bArray[2][20] ), 
        .D(\bArray[3][20] ), .S0(n7206), .S1(n7218), .Y(n7027) );
  OA22XL U9636 ( .A0(\xArray[5][23] ), .A1(n8195), .B0(\xArray[1][23] ), .B1(
        n8269), .Y(n906) );
  OA22XL U9637 ( .A0(\xArray[5][24] ), .A1(n8195), .B0(\xArray[1][24] ), .B1(
        n8269), .Y(n903) );
  AOI2BB2XL U9638 ( .B0(n9206), .B1(n8210), .A0N(\xArray[10][24] ), .A1N(n8259), .Y(n2104) );
  AOI2BB2XL U9639 ( .B0(n9198), .B1(n8210), .A0N(\xArray[10][25] ), .A1N(n8257), .Y(n2095) );
  OA22XL U9640 ( .A0(\xArray[0][27] ), .A1(n8192), .B0(\xArray[12][27] ), .B1(
        n8266), .Y(n2080) );
  OA22XL U9641 ( .A0(\xArray[0][26] ), .A1(n8191), .B0(\xArray[12][26] ), .B1(
        n8267), .Y(n2089) );
  AOI2BB2XL U9642 ( .B0(n9200), .B1(n8207), .A0N(\xArray[15][24] ), .A1N(n8255), .Y(n1174) );
  AOI2BB2XL U9643 ( .B0(n9208), .B1(n8208), .A0N(\xArray[15][23] ), .A1N(n8255), .Y(n1179) );
  OA22XL U9644 ( .A0(\xArray[4][24] ), .A1(n8197), .B0(\xArray[0][24] ), .B1(
        n8267), .Y(n1173) );
  OA22XL U9645 ( .A0(\xArray[15][27] ), .A1(n8192), .B0(\xArray[11][27] ), 
        .B1(n8266), .Y(n2079) );
  OA22XL U9646 ( .A0(\xArray[15][26] ), .A1(n8191), .B0(\xArray[11][26] ), 
        .B1(n8267), .Y(n2088) );
  OA22XL U9647 ( .A0(\xArray[1][26] ), .A1(n8188), .B0(\xArray[13][26] ), .B1(
        n8261), .Y(n1665) );
  OA22XL U9648 ( .A0(\xArray[1][25] ), .A1(n8188), .B0(\xArray[13][25] ), .B1(
        n8261), .Y(n1668) );
  AOI22XL U9649 ( .A0(n8058), .A1(n7431), .B0(\xArray[8][28] ), .B1(n8056), 
        .Y(n3189) );
  AOI22XL U9650 ( .A0(n2599), .A1(n7431), .B0(\xArray[2][28] ), .B1(n8134), 
        .Y(n2670) );
  AOI22XL U9651 ( .A0(n8058), .A1(n7429), .B0(\xArray[8][27] ), .B1(n8057), 
        .Y(n3190) );
  AOI22XL U9652 ( .A0(n8135), .A1(n7429), .B0(\xArray[2][27] ), .B1(n2601), 
        .Y(n2672) );
  OA22XL U9653 ( .A0(n8322), .A1(n1478), .B0(n7729), .B1(n1688), .Y(n2153) );
  OA22XL U9654 ( .A0(n8322), .A1(n1474), .B0(n7729), .B1(n1685), .Y(n2144) );
  MX4XL U9655 ( .A(\bArray[4][21] ), .B(\bArray[5][21] ), .C(\bArray[6][21] ), 
        .D(\bArray[7][21] ), .S0(n7206), .S1(n7218), .Y(n7030) );
  MX4XL U9656 ( .A(\bArray[12][21] ), .B(\bArray[13][21] ), .C(
        \bArray[14][21] ), .D(\bArray[15][21] ), .S0(n7206), .S1(n7218), .Y(
        n7028) );
  MX4XL U9657 ( .A(\bArray[8][21] ), .B(\bArray[9][21] ), .C(\bArray[10][21] ), 
        .D(\bArray[11][21] ), .S0(n7206), .S1(n7218), .Y(n7029) );
  INVXL U9658 ( .A(\xArray[14][21] ), .Y(n9230) );
  INVXL U9659 ( .A(\xArray[14][22] ), .Y(n9222) );
  INVXL U9660 ( .A(\xArray[5][12] ), .Y(n9298) );
  INVXL U9661 ( .A(\xArray[5][13] ), .Y(n9290) );
  INVXL U9662 ( .A(\xArray[3][20] ), .Y(n9232) );
  INVXL U9663 ( .A(\xArray[3][21] ), .Y(n9224) );
  INVXL U9664 ( .A(\xArray[9][12] ), .Y(n9300) );
  INVXL U9665 ( .A(\xArray[9][13] ), .Y(n9292) );
  INVXL U9666 ( .A(\xArray[6][11] ), .Y(n9307) );
  INVXL U9667 ( .A(\xArray[6][12] ), .Y(n9299) );
  INVXL U9668 ( .A(\xArray[10][11] ), .Y(n9309) );
  INVXL U9669 ( .A(\xArray[10][12] ), .Y(n9301) );
  MX4XL U9670 ( .A(\bArray[0][22] ), .B(\bArray[1][22] ), .C(\bArray[2][22] ), 
        .D(\bArray[3][22] ), .S0(n7207), .S1(n7219), .Y(n7035) );
  OA22XL U9671 ( .A0(\xArray[5][25] ), .A1(n8195), .B0(\xArray[1][25] ), .B1(
        n8269), .Y(n900) );
  AOI2BB2XL U9672 ( .B0(n9182), .B1(n8217), .A0N(\xArray[10][27] ), .A1N(n8257), .Y(n2077) );
  AOI2BB2XL U9673 ( .B0(n9190), .B1(n8210), .A0N(\xArray[10][26] ), .A1N(n8257), .Y(n2086) );
  OA22XL U9674 ( .A0(\xArray[0][28] ), .A1(n8192), .B0(\xArray[12][28] ), .B1(
        n8266), .Y(n2071) );
  OA22XL U9675 ( .A0(\xArray[14][27] ), .A1(n8272), .B0(\xArray[2][27] ), .B1(
        n8185), .Y(n1443) );
  OA22XL U9676 ( .A0(\xArray[4][25] ), .A1(n8197), .B0(\xArray[0][25] ), .B1(
        n8267), .Y(n1168) );
  OA22XL U9677 ( .A0(\xArray[15][28] ), .A1(n8192), .B0(\xArray[11][28] ), 
        .B1(n8266), .Y(n2070) );
  OA22XL U9678 ( .A0(\xArray[1][27] ), .A1(n8188), .B0(\xArray[13][27] ), .B1(
        n8262), .Y(n1662) );
  AOI22XL U9679 ( .A0(n3153), .A1(n7427), .B0(\xArray[8][26] ), .B1(n8057), 
        .Y(n3191) );
  AOI22XL U9680 ( .A0(n8136), .A1(n7427), .B0(\xArray[2][26] ), .B1(n2601), 
        .Y(n2674) );
  AOI22XL U9681 ( .A0(n3153), .A1(n7425), .B0(\xArray[8][25] ), .B1(n8057), 
        .Y(n3192) );
  AOI22XL U9682 ( .A0(n8135), .A1(n7425), .B0(\xArray[2][25] ), .B1(n2601), 
        .Y(n2676) );
  AOI22XL U9683 ( .A0(n8058), .A1(n7423), .B0(\xArray[8][24] ), .B1(n8057), 
        .Y(n3193) );
  AOI22XL U9684 ( .A0(n8136), .A1(n7423), .B0(\xArray[2][24] ), .B1(n2601), 
        .Y(n2678) );
  OA22XL U9685 ( .A0(n8322), .A1(n1470), .B0(n7729), .B1(n1682), .Y(n2135) );
  MX4XL U9686 ( .A(\bArray[4][23] ), .B(\bArray[5][23] ), .C(\bArray[6][23] ), 
        .D(\bArray[7][23] ), .S0(n7207), .S1(n7219), .Y(n7038) );
  MX4XL U9687 ( .A(\bArray[12][23] ), .B(\bArray[13][23] ), .C(
        \bArray[14][23] ), .D(\bArray[15][23] ), .S0(n7207), .S1(n7219), .Y(
        n7036) );
  MX4XL U9688 ( .A(\bArray[8][23] ), .B(\bArray[9][23] ), .C(\bArray[10][23] ), 
        .D(\bArray[11][23] ), .S0(n7207), .S1(n7219), .Y(n7037) );
  MX4XL U9689 ( .A(\bArray[4][24] ), .B(\bArray[5][24] ), .C(\bArray[6][24] ), 
        .D(\bArray[7][24] ), .S0(n7207), .S1(n7219), .Y(n7042) );
  MX4XL U9690 ( .A(\bArray[12][24] ), .B(\bArray[13][24] ), .C(
        \bArray[14][24] ), .D(\bArray[15][24] ), .S0(n7207), .S1(n7219), .Y(
        n7040) );
  MX4XL U9691 ( .A(\bArray[8][24] ), .B(\bArray[9][24] ), .C(\bArray[10][24] ), 
        .D(\bArray[11][24] ), .S0(n7207), .S1(n7219), .Y(n7041) );
  INVXL U9692 ( .A(\xArray[14][23] ), .Y(n9214) );
  INVXL U9693 ( .A(\xArray[14][24] ), .Y(n9206) );
  INVXL U9694 ( .A(\xArray[5][14] ), .Y(n9282) );
  INVXL U9695 ( .A(\xArray[5][15] ), .Y(n9274) );
  AOI2BB2XL U9696 ( .B0(n9192), .B1(n8217), .A0N(\xArray[15][25] ), .A1N(n8255), .Y(n1169) );
  INVXL U9697 ( .A(\xArray[3][22] ), .Y(n9216) );
  INVXL U9698 ( .A(\xArray[3][23] ), .Y(n9208) );
  INVXL U9699 ( .A(\xArray[9][14] ), .Y(n9284) );
  INVXL U9700 ( .A(\xArray[9][15] ), .Y(n9276) );
  INVXL U9701 ( .A(\xArray[6][13] ), .Y(n9291) );
  INVXL U9702 ( .A(\xArray[6][14] ), .Y(n9283) );
  INVXL U9703 ( .A(\xArray[10][13] ), .Y(n9293) );
  INVXL U9704 ( .A(\xArray[10][14] ), .Y(n9285) );
  MX4XL U9705 ( .A(\bArray[0][23] ), .B(\bArray[1][23] ), .C(\bArray[2][23] ), 
        .D(\bArray[3][23] ), .S0(n7207), .S1(n7219), .Y(n7039) );
  MX4XL U9706 ( .A(\bArray[0][24] ), .B(\bArray[1][24] ), .C(\bArray[2][24] ), 
        .D(\bArray[3][24] ), .S0(n7207), .S1(n7219), .Y(n7043) );
  OA22XL U9707 ( .A0(\xArray[5][27] ), .A1(n8195), .B0(\xArray[1][27] ), .B1(
        n8269), .Y(n894) );
  OA22XL U9708 ( .A0(\xArray[5][26] ), .A1(n8195), .B0(\xArray[1][26] ), .B1(
        n8269), .Y(n897) );
  AOI2BB2XL U9709 ( .B0(n9166), .B1(n8203), .A0N(\xArray[10][29] ), .A1N(n8256), .Y(n2059) );
  OA22XL U9710 ( .A0(\xArray[0][30] ), .A1(n8192), .B0(\xArray[12][30] ), .B1(
        n8266), .Y(n2053) );
  AOI2BB2XL U9711 ( .B0(n9168), .B1(n8212), .A0N(\xArray[15][28] ), .A1N(n8256), .Y(n1154) );
  OA22XL U9712 ( .A0(\xArray[4][28] ), .A1(n8197), .B0(\xArray[0][28] ), .B1(
        n8267), .Y(n1153) );
  OA22XL U9713 ( .A0(\xArray[14][30] ), .A1(n8271), .B0(\xArray[2][30] ), .B1(
        n8185), .Y(n1431) );
  OA22XL U9714 ( .A0(\xArray[15][30] ), .A1(n8192), .B0(\xArray[11][30] ), 
        .B1(n8266), .Y(n2052) );
  OA22XL U9715 ( .A0(\xArray[1][30] ), .A1(n8189), .B0(\xArray[13][30] ), .B1(
        n8266), .Y(n1653) );
  AOI22XL U9716 ( .A0(n8058), .A1(n7421), .B0(\xArray[8][23] ), .B1(n8057), 
        .Y(n3194) );
  AOI22XL U9717 ( .A0(n8135), .A1(n7421), .B0(\xArray[2][23] ), .B1(n2601), 
        .Y(n2680) );
  AOI22XL U9718 ( .A0(n8058), .A1(n7419), .B0(\xArray[8][22] ), .B1(n8057), 
        .Y(n3195) );
  AOI22XL U9719 ( .A0(n8136), .A1(n7419), .B0(\xArray[2][22] ), .B1(n2601), 
        .Y(n2682) );
  AOI22XL U9720 ( .A0(n8058), .A1(n7417), .B0(\xArray[8][21] ), .B1(n8057), 
        .Y(n3196) );
  AOI22XL U9721 ( .A0(n8136), .A1(n7417), .B0(\xArray[2][21] ), .B1(n2601), 
        .Y(n2684) );
  OAI22XL U9722 ( .A0(\xArray[10][22] ), .A1(n7892), .B0(n7898), .B1(n7419), 
        .Y(n3338) );
  OAI22XL U9723 ( .A0(\xArray[13][22] ), .A1(n7869), .B0(n7882), .B1(n7419), 
        .Y(n3543) );
  OAI22XL U9724 ( .A0(\xArray[10][21] ), .A1(n7892), .B0(n7898), .B1(n7417), 
        .Y(n3339) );
  OAI22XL U9725 ( .A0(\xArray[13][21] ), .A1(n7869), .B0(n7882), .B1(n7417), 
        .Y(n3544) );
  OAI22XL U9726 ( .A0(\xArray[1][23] ), .A1(n7790), .B0(n7801), .B1(n7421), 
        .Y(n2570) );
  OAI22XL U9727 ( .A0(\xArray[10][23] ), .A1(n7892), .B0(n7899), .B1(n7421), 
        .Y(n3337) );
  OAI22XL U9728 ( .A0(\xArray[13][23] ), .A1(n7869), .B0(n7882), .B1(n7421), 
        .Y(n3542) );
  OAI22XL U9729 ( .A0(\xArray[1][22] ), .A1(n7790), .B0(n7802), .B1(n7419), 
        .Y(n2571) );
  OAI22XL U9730 ( .A0(\xArray[1][21] ), .A1(n7789), .B0(n7802), .B1(n7417), 
        .Y(n2572) );
  OAI22XL U9731 ( .A0(\xArray[0][23] ), .A1(n7769), .B0(n7777), .B1(n7421), 
        .Y(n2452) );
  OAI22XL U9732 ( .A0(\xArray[0][22] ), .A1(n7769), .B0(n7777), .B1(n7419), 
        .Y(n2455) );
  OAI22XL U9733 ( .A0(\xArray[0][21] ), .A1(n7769), .B0(n7778), .B1(n7417), 
        .Y(n2458) );
  OAI22XL U9734 ( .A0(\xArray[11][23] ), .A1(n7830), .B0(n7844), .B1(n7421), 
        .Y(n3405) );
  OAI22XL U9735 ( .A0(\xArray[11][22] ), .A1(n7830), .B0(n7838), .B1(n7419), 
        .Y(n3406) );
  OAI22XL U9736 ( .A0(\xArray[11][21] ), .A1(n7830), .B0(n7838), .B1(n7417), 
        .Y(n3407) );
  OAI22XL U9737 ( .A0(\xArray[6][22] ), .A1(n7810), .B0(n7818), .B1(n7419), 
        .Y(n3054) );
  OAI22XL U9738 ( .A0(\xArray[6][21] ), .A1(n7810), .B0(n7818), .B1(n7417), 
        .Y(n3055) );
  OAI22XL U9739 ( .A0(\xArray[7][23] ), .A1(n7849), .B0(n7858), .B1(n7421), 
        .Y(n3124) );
  OAI22XL U9740 ( .A0(\xArray[12][23] ), .A1(n7912), .B0(n7919), .B1(n7421), 
        .Y(n3474) );
  OAI22XL U9741 ( .A0(\xArray[7][22] ), .A1(n7849), .B0(n7857), .B1(n7419), 
        .Y(n3125) );
  OAI22XL U9742 ( .A0(\xArray[12][22] ), .A1(n7912), .B0(n7918), .B1(n7419), 
        .Y(n3475) );
  OAI22XL U9743 ( .A0(\xArray[7][21] ), .A1(n7849), .B0(n7857), .B1(n7417), 
        .Y(n3126) );
  OAI22XL U9744 ( .A0(\xArray[12][21] ), .A1(n7912), .B0(n7918), .B1(n7417), 
        .Y(n3476) );
  OA22XL U9745 ( .A0(n8322), .A1(n1466), .B0(n7729), .B1(n1679), .Y(n2126) );
  MX4XL U9746 ( .A(\bArray[4][26] ), .B(\bArray[5][26] ), .C(\bArray[6][26] ), 
        .D(\bArray[7][26] ), .S0(n7208), .S1(n7220), .Y(n7050) );
  MX4XL U9747 ( .A(\bArray[12][26] ), .B(\bArray[13][26] ), .C(
        \bArray[14][26] ), .D(\bArray[15][26] ), .S0(n7208), .S1(n7220), .Y(
        n7048) );
  MX4XL U9748 ( .A(\bArray[8][26] ), .B(\bArray[9][26] ), .C(\bArray[10][26] ), 
        .D(\bArray[11][26] ), .S0(n7208), .S1(n7220), .Y(n7049) );
  INVXL U9749 ( .A(\xArray[14][25] ), .Y(n9198) );
  INVXL U9750 ( .A(\xArray[14][26] ), .Y(n9190) );
  INVXL U9751 ( .A(\xArray[5][16] ), .Y(n9266) );
  INVXL U9752 ( .A(\xArray[5][17] ), .Y(n9258) );
  INVXL U9753 ( .A(\xArray[3][24] ), .Y(n9200) );
  INVXL U9754 ( .A(\xArray[3][25] ), .Y(n9192) );
  INVXL U9755 ( .A(\xArray[9][16] ), .Y(n9268) );
  INVXL U9756 ( .A(\xArray[9][17] ), .Y(n9260) );
  INVXL U9757 ( .A(\xArray[6][15] ), .Y(n9275) );
  INVXL U9758 ( .A(\xArray[6][16] ), .Y(n9267) );
  INVXL U9759 ( .A(\xArray[10][15] ), .Y(n9277) );
  INVXL U9760 ( .A(\xArray[10][16] ), .Y(n9269) );
  MX4XL U9761 ( .A(\bArray[0][26] ), .B(\bArray[1][26] ), .C(\bArray[2][26] ), 
        .D(\bArray[3][26] ), .S0(n7208), .S1(n7220), .Y(n7051) );
  OA22XL U9762 ( .A0(\xArray[5][28] ), .A1(n8195), .B0(\xArray[1][28] ), .B1(
        n8269), .Y(n891) );
  AOI2BB2XL U9763 ( .B0(n9150), .B1(n8203), .A0N(\xArray[10][31] ), .A1N(n8256), .Y(n2041) );
  AOI2BB2XL U9764 ( .B0(n9158), .B1(n6693), .A0N(\xArray[10][30] ), .A1N(n8256), .Y(n2050) );
  AOI2BB2XL U9765 ( .B0(n9152), .B1(n8212), .A0N(\xArray[15][30] ), .A1N(n8256), .Y(n1144) );
  OA22XL U9766 ( .A0(\xArray[4][29] ), .A1(n8197), .B0(\xArray[0][29] ), .B1(
        n8267), .Y(n1148) );
  OA22XL U9767 ( .A0(\xArray[4][30] ), .A1(n8197), .B0(\xArray[0][30] ), .B1(
        n8267), .Y(n1143) );
  OA22XL U9768 ( .A0(\xArray[14][31] ), .A1(n8271), .B0(\xArray[2][31] ), .B1(
        n8185), .Y(n1427) );
  OA22XL U9769 ( .A0(\xArray[15][31] ), .A1(n8192), .B0(\xArray[11][31] ), 
        .B1(n8266), .Y(n2043) );
  OA22XL U9770 ( .A0(\xArray[15][32] ), .A1(n8192), .B0(\xArray[11][32] ), 
        .B1(n8266), .Y(n2034) );
  OA22XL U9771 ( .A0(\xArray[1][31] ), .A1(n8200), .B0(\xArray[13][31] ), .B1(
        n8270), .Y(n1650) );
  AOI22XL U9772 ( .A0(n8058), .A1(n7415), .B0(\xArray[8][20] ), .B1(n8057), 
        .Y(n3197) );
  AOI22XL U9773 ( .A0(n8136), .A1(n7415), .B0(\xArray[2][20] ), .B1(n2601), 
        .Y(n2686) );
  AOI22XL U9774 ( .A0(n8058), .A1(n7413), .B0(\xArray[8][19] ), .B1(n8057), 
        .Y(n3198) );
  AOI22XL U9775 ( .A0(n8137), .A1(n7413), .B0(\xArray[2][19] ), .B1(n2601), 
        .Y(n2688) );
  AOI22XL U9776 ( .A0(n8060), .A1(n7411), .B0(\xArray[8][18] ), .B1(n8057), 
        .Y(n3199) );
  AOI22XL U9777 ( .A0(n8135), .A1(n7411), .B0(\xArray[2][18] ), .B1(n2601), 
        .Y(n2690) );
  OAI22XL U9778 ( .A0(\xArray[1][20] ), .A1(n7790), .B0(n7802), .B1(n7415), 
        .Y(n2573) );
  OAI22XL U9779 ( .A0(\xArray[10][20] ), .A1(n7892), .B0(n7898), .B1(n7415), 
        .Y(n3340) );
  OAI22XL U9780 ( .A0(\xArray[13][20] ), .A1(n7869), .B0(n7882), .B1(n7415), 
        .Y(n3545) );
  OAI22XL U9781 ( .A0(\xArray[1][19] ), .A1(n7790), .B0(n7802), .B1(n7413), 
        .Y(n2574) );
  OAI22XL U9782 ( .A0(\xArray[10][19] ), .A1(n7892), .B0(n7898), .B1(n7413), 
        .Y(n3341) );
  OAI22XL U9783 ( .A0(\xArray[13][19] ), .A1(n7869), .B0(n7882), .B1(n7413), 
        .Y(n3546) );
  OAI22XL U9784 ( .A0(\xArray[1][18] ), .A1(n7789), .B0(n7802), .B1(n7411), 
        .Y(n2575) );
  OAI22XL U9785 ( .A0(\xArray[10][18] ), .A1(n7892), .B0(n7897), .B1(n7411), 
        .Y(n3342) );
  OAI22XL U9786 ( .A0(\xArray[13][18] ), .A1(n7869), .B0(n7882), .B1(n7411), 
        .Y(n3547) );
  OAI22XL U9787 ( .A0(\xArray[0][20] ), .A1(n7769), .B0(n7778), .B1(n7415), 
        .Y(n2461) );
  OAI22XL U9788 ( .A0(\xArray[0][19] ), .A1(n7769), .B0(n7778), .B1(n7413), 
        .Y(n2464) );
  OAI22XL U9789 ( .A0(\xArray[0][18] ), .A1(n7769), .B0(n7777), .B1(n7411), 
        .Y(n2467) );
  OAI22XL U9790 ( .A0(\xArray[11][20] ), .A1(n7830), .B0(n7838), .B1(n7415), 
        .Y(n3408) );
  OAI22XL U9791 ( .A0(\xArray[11][19] ), .A1(n7830), .B0(n7838), .B1(n7413), 
        .Y(n3409) );
  OAI22XL U9792 ( .A0(\xArray[11][18] ), .A1(n7830), .B0(n7837), .B1(n7411), 
        .Y(n3410) );
  OAI22XL U9793 ( .A0(\xArray[6][20] ), .A1(n7810), .B0(n7818), .B1(n7415), 
        .Y(n3056) );
  OAI22XL U9794 ( .A0(\xArray[6][19] ), .A1(n7810), .B0(n7818), .B1(n7413), 
        .Y(n3057) );
  OAI22XL U9795 ( .A0(\xArray[6][18] ), .A1(n7810), .B0(n7817), .B1(n7411), 
        .Y(n3058) );
  OAI22XL U9796 ( .A0(\xArray[7][20] ), .A1(n7849), .B0(n7857), .B1(n7415), 
        .Y(n3127) );
  OAI22XL U9797 ( .A0(\xArray[12][20] ), .A1(n7912), .B0(n7918), .B1(n7415), 
        .Y(n3477) );
  OAI22XL U9798 ( .A0(\xArray[7][19] ), .A1(n7849), .B0(n7857), .B1(n7413), 
        .Y(n3128) );
  OAI22XL U9799 ( .A0(\xArray[12][19] ), .A1(n7912), .B0(n7918), .B1(n7413), 
        .Y(n3478) );
  OAI22XL U9800 ( .A0(\xArray[7][18] ), .A1(n7849), .B0(n7856), .B1(n7411), 
        .Y(n3129) );
  OAI22XL U9801 ( .A0(\xArray[12][18] ), .A1(n7912), .B0(n7917), .B1(n7411), 
        .Y(n3479) );
  MX4XL U9802 ( .A(\bArray[4][27] ), .B(\bArray[5][27] ), .C(\bArray[6][27] ), 
        .D(\bArray[7][27] ), .S0(n7208), .S1(n7220), .Y(n7054) );
  MX4XL U9803 ( .A(\bArray[12][27] ), .B(\bArray[13][27] ), .C(
        \bArray[14][27] ), .D(\bArray[15][27] ), .S0(n7208), .S1(n7220), .Y(
        n7052) );
  MX4XL U9804 ( .A(\bArray[8][27] ), .B(\bArray[9][27] ), .C(\bArray[10][27] ), 
        .D(\bArray[11][27] ), .S0(n7208), .S1(n7220), .Y(n7053) );
  MX4XL U9805 ( .A(\bArray[12][28] ), .B(\bArray[13][28] ), .C(
        \bArray[14][28] ), .D(\bArray[15][28] ), .S0(n7208), .S1(n7220), .Y(
        n7056) );
  INVXL U9806 ( .A(\xArray[14][27] ), .Y(n9182) );
  INVXL U9807 ( .A(\xArray[14][28] ), .Y(n9174) );
  INVXL U9808 ( .A(\xArray[5][18] ), .Y(n9250) );
  INVXL U9809 ( .A(\xArray[5][19] ), .Y(n9242) );
  AOI2BB2XL U9810 ( .B0(n9160), .B1(n8212), .A0N(\xArray[15][29] ), .A1N(n8256), .Y(n1149) );
  INVXL U9811 ( .A(\xArray[3][26] ), .Y(n9184) );
  INVXL U9812 ( .A(\xArray[3][27] ), .Y(n9176) );
  INVXL U9813 ( .A(\xArray[9][18] ), .Y(n9252) );
  INVXL U9814 ( .A(\xArray[9][19] ), .Y(n9244) );
  INVXL U9815 ( .A(\xArray[6][17] ), .Y(n9259) );
  INVXL U9816 ( .A(\xArray[6][18] ), .Y(n9251) );
  INVXL U9817 ( .A(\xArray[10][17] ), .Y(n9261) );
  INVXL U9818 ( .A(\xArray[10][18] ), .Y(n9253) );
  MX4XL U9819 ( .A(\bArray[0][27] ), .B(\bArray[1][27] ), .C(\bArray[2][27] ), 
        .D(\bArray[3][27] ), .S0(n7208), .S1(n7220), .Y(n7055) );
  OA22XL U9820 ( .A0(\xArray[14][32] ), .A1(n8271), .B0(\xArray[2][32] ), .B1(
        n8185), .Y(n1423) );
  OA22XL U9821 ( .A0(\xArray[0][31] ), .A1(n8192), .B0(\xArray[12][31] ), .B1(
        n8266), .Y(n2044) );
  OA22XL U9822 ( .A0(\xArray[0][32] ), .A1(n8192), .B0(\xArray[12][32] ), .B1(
        n8266), .Y(n2035) );
  OA22XL U9823 ( .A0(\xArray[5][29] ), .A1(n8195), .B0(\xArray[1][29] ), .B1(
        n8269), .Y(n888) );
  AOI2BB2XL U9824 ( .B0(n9142), .B1(n8214), .A0N(\xArray[10][32] ), .A1N(n8256), .Y(n2032) );
  OA22XL U9825 ( .A0(\xArray[5][31] ), .A1(n8195), .B0(\xArray[1][31] ), .B1(
        n8267), .Y(n882) );
  AOI2BB2XL U9826 ( .B0(n9134), .B1(n8203), .A0N(\xArray[10][33] ), .A1N(n8255), .Y(n2023) );
  OA22XL U9827 ( .A0(\xArray[0][34] ), .A1(n8192), .B0(\xArray[12][34] ), .B1(
        n8265), .Y(n2017) );
  AOI2BB2XL U9828 ( .B0(n9144), .B1(n8212), .A0N(\xArray[15][31] ), .A1N(n8256), .Y(n1139) );
  OA22XL U9829 ( .A0(\xArray[14][34] ), .A1(n8271), .B0(\xArray[2][34] ), .B1(
        n8185), .Y(n1415) );
  OA22XL U9830 ( .A0(\xArray[15][33] ), .A1(n8192), .B0(\xArray[11][33] ), 
        .B1(n8265), .Y(n2025) );
  OA22XL U9831 ( .A0(\xArray[15][34] ), .A1(n8192), .B0(\xArray[11][34] ), 
        .B1(n8265), .Y(n2016) );
  AOI22XL U9832 ( .A0(n8060), .A1(n7409), .B0(\xArray[8][17] ), .B1(n8057), 
        .Y(n3200) );
  AOI22XL U9833 ( .A0(n8136), .A1(n7409), .B0(\xArray[2][17] ), .B1(n8134), 
        .Y(n2692) );
  AOI22XL U9834 ( .A0(n8059), .A1(n7407), .B0(\xArray[8][16] ), .B1(n8057), 
        .Y(n3201) );
  AOI22XL U9835 ( .A0(n8137), .A1(n7407), .B0(\xArray[2][16] ), .B1(n8132), 
        .Y(n2694) );
  AOI22XL U9836 ( .A0(n8060), .A1(n7405), .B0(\xArray[8][15] ), .B1(n3154), 
        .Y(n3202) );
  AOI22XL U9837 ( .A0(n8137), .A1(n7405), .B0(\xArray[2][15] ), .B1(n8134), 
        .Y(n2696) );
  OAI22XL U9838 ( .A0(\xArray[1][17] ), .A1(n7789), .B0(n7800), .B1(n7409), 
        .Y(n2576) );
  OAI22XL U9839 ( .A0(\xArray[10][17] ), .A1(n7892), .B0(n7897), .B1(n7409), 
        .Y(n3343) );
  OAI22XL U9840 ( .A0(\xArray[13][17] ), .A1(n7869), .B0(n7882), .B1(n7409), 
        .Y(n3548) );
  OAI22XL U9841 ( .A0(\xArray[1][16] ), .A1(n7788), .B0(n7802), .B1(n7407), 
        .Y(n2577) );
  OAI22XL U9842 ( .A0(\xArray[10][16] ), .A1(n7892), .B0(n7897), .B1(n7407), 
        .Y(n3344) );
  OAI22XL U9843 ( .A0(\xArray[13][16] ), .A1(n7869), .B0(n7882), .B1(n7407), 
        .Y(n3549) );
  OAI22XL U9844 ( .A0(\xArray[1][15] ), .A1(n7788), .B0(n7801), .B1(n7405), 
        .Y(n2578) );
  OAI22XL U9845 ( .A0(\xArray[10][15] ), .A1(n7893), .B0(n7897), .B1(n7405), 
        .Y(n3345) );
  OAI22XL U9846 ( .A0(\xArray[13][15] ), .A1(n7870), .B0(n7880), .B1(n7405), 
        .Y(n3550) );
  OAI22XL U9847 ( .A0(\xArray[0][17] ), .A1(n7769), .B0(n7778), .B1(n7409), 
        .Y(n2470) );
  OAI22XL U9848 ( .A0(\xArray[0][16] ), .A1(n7769), .B0(n7777), .B1(n7407), 
        .Y(n2473) );
  OAI22XL U9849 ( .A0(\xArray[0][15] ), .A1(n7770), .B0(n7778), .B1(n7405), 
        .Y(n2476) );
  OAI22XL U9850 ( .A0(\xArray[11][17] ), .A1(n7830), .B0(n7837), .B1(n7409), 
        .Y(n3411) );
  OAI22XL U9851 ( .A0(\xArray[11][16] ), .A1(n7830), .B0(n7837), .B1(n7407), 
        .Y(n3412) );
  OAI22XL U9852 ( .A0(\xArray[11][15] ), .A1(n7831), .B0(n7837), .B1(n7405), 
        .Y(n3413) );
  OAI22XL U9853 ( .A0(\xArray[6][17] ), .A1(n7810), .B0(n7817), .B1(n7409), 
        .Y(n3059) );
  OAI22XL U9854 ( .A0(\xArray[6][16] ), .A1(n7810), .B0(n7817), .B1(n7407), 
        .Y(n3060) );
  OAI22XL U9855 ( .A0(\xArray[6][15] ), .A1(n7811), .B0(n7817), .B1(n7405), 
        .Y(n3061) );
  OAI22XL U9856 ( .A0(\xArray[7][17] ), .A1(n7849), .B0(n7856), .B1(n7409), 
        .Y(n3130) );
  OAI22XL U9857 ( .A0(\xArray[12][17] ), .A1(n7912), .B0(n7917), .B1(n7409), 
        .Y(n3480) );
  OAI22XL U9858 ( .A0(\xArray[7][16] ), .A1(n7849), .B0(n7856), .B1(n7407), 
        .Y(n3131) );
  OAI22XL U9859 ( .A0(\xArray[12][16] ), .A1(n7912), .B0(n7917), .B1(n7407), 
        .Y(n3481) );
  OAI22XL U9860 ( .A0(\xArray[7][15] ), .A1(n7850), .B0(n7856), .B1(n7405), 
        .Y(n3132) );
  OAI22XL U9861 ( .A0(\xArray[12][15] ), .A1(n7913), .B0(n7917), .B1(n7405), 
        .Y(n3482) );
  MX4XL U9862 ( .A(\bArray[4][29] ), .B(\bArray[5][29] ), .C(\bArray[6][29] ), 
        .D(\bArray[7][29] ), .S0(n7209), .S1(n7221), .Y(n7062) );
  MX4XL U9863 ( .A(\bArray[12][29] ), .B(\bArray[13][29] ), .C(
        \bArray[14][29] ), .D(\bArray[15][29] ), .S0(n7209), .S1(n7221), .Y(
        n7060) );
  MX4XL U9864 ( .A(\bArray[8][29] ), .B(\bArray[9][29] ), .C(\bArray[10][29] ), 
        .D(\bArray[11][29] ), .S0(n7209), .S1(n7221), .Y(n7061) );
  MX4XL U9865 ( .A(\bArray[4][30] ), .B(\bArray[5][30] ), .C(\bArray[6][30] ), 
        .D(\bArray[7][30] ), .S0(n7209), .S1(n7221), .Y(n7066) );
  MX4XL U9866 ( .A(\bArray[12][30] ), .B(\bArray[13][30] ), .C(
        \bArray[14][30] ), .D(\bArray[15][30] ), .S0(n7209), .S1(n7221), .Y(
        n7064) );
  MX4XL U9867 ( .A(\bArray[8][30] ), .B(\bArray[9][30] ), .C(\bArray[10][30] ), 
        .D(\bArray[11][30] ), .S0(n7209), .S1(n7221), .Y(n7065) );
  INVXL U9868 ( .A(\xArray[14][29] ), .Y(n9166) );
  INVXL U9869 ( .A(\xArray[14][30] ), .Y(n9158) );
  INVXL U9870 ( .A(\xArray[5][20] ), .Y(n9234) );
  INVXL U9871 ( .A(\xArray[5][21] ), .Y(n9226) );
  INVXL U9872 ( .A(\xArray[3][28] ), .Y(n9168) );
  INVXL U9873 ( .A(\xArray[3][29] ), .Y(n9160) );
  INVXL U9874 ( .A(\xArray[9][20] ), .Y(n9236) );
  INVXL U9875 ( .A(\xArray[9][21] ), .Y(n9228) );
  INVXL U9876 ( .A(\xArray[6][19] ), .Y(n9243) );
  INVXL U9877 ( .A(\xArray[6][20] ), .Y(n9235) );
  INVXL U9878 ( .A(\xArray[10][19] ), .Y(n9245) );
  INVXL U9879 ( .A(\xArray[10][20] ), .Y(n9237) );
  MX4XL U9880 ( .A(\bArray[0][29] ), .B(\bArray[1][29] ), .C(\bArray[2][29] ), 
        .D(\bArray[3][29] ), .S0(n7209), .S1(n7221), .Y(n7063) );
  MX4XL U9881 ( .A(\bArray[0][30] ), .B(\bArray[1][30] ), .C(\bArray[2][30] ), 
        .D(\bArray[3][30] ), .S0(n7209), .S1(n7221), .Y(n7067) );
  OA22XL U9882 ( .A0(\xArray[14][33] ), .A1(n8272), .B0(\xArray[2][33] ), .B1(
        n8185), .Y(n1419) );
  OA22XL U9883 ( .A0(\xArray[0][33] ), .A1(n8192), .B0(\xArray[12][33] ), .B1(
        n8265), .Y(n2026) );
  OA22XL U9884 ( .A0(\xArray[5][30] ), .A1(n8195), .B0(\xArray[1][30] ), .B1(
        n8269), .Y(n885) );
  OA22XL U9885 ( .A0(\xArray[5][32] ), .A1(n8195), .B0(\xArray[1][32] ), .B1(
        n8267), .Y(n879) );
  AOI2BB2XL U9886 ( .B0(n9118), .B1(n8217), .A0N(\xArray[10][35] ), .A1N(n8255), .Y(n2005) );
  AOI2BB2XL U9887 ( .B0(n9128), .B1(n8217), .A0N(\xArray[15][33] ), .A1N(n8256), .Y(n1129) );
  AOI2BB2XL U9888 ( .B0(n9120), .B1(n8217), .A0N(\xArray[15][34] ), .A1N(n8256), .Y(n1124) );
  OA22XL U9889 ( .A0(\xArray[14][35] ), .A1(n8271), .B0(\xArray[2][35] ), .B1(
        n8185), .Y(n1411) );
  AOI22XL U9890 ( .A0(n8060), .A1(n7403), .B0(\xArray[8][14] ), .B1(n3154), 
        .Y(n3203) );
  AOI22XL U9891 ( .A0(n8137), .A1(n7403), .B0(\xArray[2][14] ), .B1(n8134), 
        .Y(n2698) );
  AOI22XL U9892 ( .A0(n8060), .A1(n7401), .B0(\xArray[8][13] ), .B1(n3154), 
        .Y(n3204) );
  AOI22XL U9893 ( .A0(n8137), .A1(n7401), .B0(\xArray[2][13] ), .B1(n8134), 
        .Y(n2700) );
  OAI22XL U9894 ( .A0(\xArray[1][14] ), .A1(n7789), .B0(n7801), .B1(n7403), 
        .Y(n2579) );
  OAI22XL U9895 ( .A0(\xArray[10][14] ), .A1(n7893), .B0(n7896), .B1(n7403), 
        .Y(n3346) );
  OAI22XL U9896 ( .A0(\xArray[13][14] ), .A1(n7869), .B0(n7880), .B1(n7403), 
        .Y(n3551) );
  OAI22XL U9897 ( .A0(\xArray[1][13] ), .A1(n7788), .B0(n7801), .B1(n7401), 
        .Y(n2580) );
  OAI22XL U9898 ( .A0(\xArray[10][13] ), .A1(n7893), .B0(n7896), .B1(n7401), 
        .Y(n3347) );
  OAI22XL U9899 ( .A0(\xArray[13][13] ), .A1(n7868), .B0(n7880), .B1(n7401), 
        .Y(n3552) );
  OAI22XL U9900 ( .A0(\xArray[0][14] ), .A1(n7769), .B0(n7777), .B1(n7403), 
        .Y(n2479) );
  OAI22XL U9901 ( .A0(\xArray[0][13] ), .A1(n7768), .B0(n7777), .B1(n7401), 
        .Y(n2482) );
  OAI22XL U9902 ( .A0(\xArray[11][14] ), .A1(n7831), .B0(n7836), .B1(n7403), 
        .Y(n3414) );
  OAI22XL U9903 ( .A0(\xArray[11][13] ), .A1(n7831), .B0(n7836), .B1(n7401), 
        .Y(n3415) );
  OAI22XL U9904 ( .A0(\xArray[11][12] ), .A1(n7831), .B0(n7836), .B1(n7399), 
        .Y(n3416) );
  OAI22XL U9905 ( .A0(\xArray[6][14] ), .A1(n7811), .B0(n7816), .B1(n7403), 
        .Y(n3062) );
  OAI22XL U9906 ( .A0(\xArray[6][13] ), .A1(n7811), .B0(n7816), .B1(n7401), 
        .Y(n3063) );
  OAI22XL U9907 ( .A0(\xArray[6][12] ), .A1(n7811), .B0(n7816), .B1(n7399), 
        .Y(n3064) );
  OAI22XL U9908 ( .A0(\xArray[7][14] ), .A1(n7850), .B0(n7855), .B1(n7403), 
        .Y(n3133) );
  OAI22XL U9909 ( .A0(\xArray[12][14] ), .A1(n7913), .B0(n7926), .B1(n7403), 
        .Y(n3483) );
  OAI22XL U9910 ( .A0(\xArray[7][13] ), .A1(n7850), .B0(n7855), .B1(n7401), 
        .Y(n3134) );
  OAI22XL U9911 ( .A0(\xArray[12][13] ), .A1(n7913), .B0(n7926), .B1(n7401), 
        .Y(n3484) );
  OAI22XL U9912 ( .A0(\xArray[7][12] ), .A1(n7850), .B0(n7855), .B1(n7399), 
        .Y(n3135) );
  OAI22XL U9913 ( .A0(\xArray[12][12] ), .A1(n7913), .B0(n7926), .B1(n7399), 
        .Y(n3485) );
  OA22XL U9914 ( .A0(n8312), .A1(n1438), .B0(n7729), .B1(n1658), .Y(n2063) );
  MX4XL U9915 ( .A(\bArray[12][31] ), .B(\bArray[13][31] ), .C(
        \bArray[14][31] ), .D(\bArray[15][31] ), .S0(n7209), .S1(n7221), .Y(
        n7068) );
  MX4XL U9916 ( .A(\bArray[8][31] ), .B(\bArray[9][31] ), .C(\bArray[10][31] ), 
        .D(\bArray[11][31] ), .S0(n7209), .S1(n7221), .Y(n7069) );
  MX4XL U9917 ( .A(\bArray[4][32] ), .B(\bArray[5][32] ), .C(\bArray[6][32] ), 
        .D(\bArray[7][32] ), .S0(n7210), .S1(n8409), .Y(n7074) );
  MX4XL U9918 ( .A(\bArray[12][32] ), .B(\bArray[13][32] ), .C(
        \bArray[14][32] ), .D(\bArray[15][32] ), .S0(n7210), .S1(n7214), .Y(
        n7072) );
  MX4XL U9919 ( .A(\bArray[8][32] ), .B(\bArray[9][32] ), .C(\bArray[10][32] ), 
        .D(\bArray[11][32] ), .S0(n7210), .S1(n8409), .Y(n7073) );
  INVXL U9920 ( .A(\xArray[14][31] ), .Y(n9150) );
  INVXL U9921 ( .A(\xArray[5][22] ), .Y(n9218) );
  INVXL U9922 ( .A(\xArray[3][30] ), .Y(n9152) );
  INVXL U9923 ( .A(\xArray[3][31] ), .Y(n9144) );
  INVXL U9924 ( .A(\xArray[9][22] ), .Y(n9220) );
  INVXL U9925 ( .A(\xArray[6][21] ), .Y(n9227) );
  INVXL U9926 ( .A(\xArray[6][22] ), .Y(n9219) );
  INVXL U9927 ( .A(\xArray[10][21] ), .Y(n9229) );
  INVXL U9928 ( .A(\xArray[10][22] ), .Y(n9221) );
  MX4XL U9929 ( .A(\bArray[0][32] ), .B(\bArray[1][32] ), .C(\bArray[2][32] ), 
        .D(\bArray[3][32] ), .S0(n7210), .S1(n8409), .Y(n7075) );
  OA22XL U9930 ( .A0(\xArray[14][36] ), .A1(n8271), .B0(\xArray[2][36] ), .B1(
        n8185), .Y(n1407) );
  OA22XL U9931 ( .A0(\xArray[4][33] ), .A1(n8197), .B0(\xArray[0][33] ), .B1(
        n8263), .Y(n1128) );
  OA22XL U9932 ( .A0(\xArray[4][34] ), .A1(n8197), .B0(\xArray[0][34] ), .B1(
        n8263), .Y(n1123) );
  OA22XL U9933 ( .A0(\xArray[0][36] ), .A1(n8192), .B0(\xArray[12][36] ), .B1(
        n8265), .Y(n1999) );
  OA22XL U9934 ( .A0(\xArray[15][36] ), .A1(n8192), .B0(\xArray[11][36] ), 
        .B1(n8265), .Y(n1998) );
  OA22XL U9935 ( .A0(\xArray[5][33] ), .A1(n8195), .B0(\xArray[1][33] ), .B1(
        n8267), .Y(n876) );
  AOI2BB2XL U9936 ( .B0(n9102), .B1(n8206), .A0N(\xArray[10][37] ), .A1N(n8255), .Y(n1987) );
  OA22XL U9937 ( .A0(\xArray[0][38] ), .A1(n8193), .B0(\xArray[12][38] ), .B1(
        n8264), .Y(n1981) );
  OA22XL U9938 ( .A0(\xArray[0][37] ), .A1(n8193), .B0(\xArray[12][37] ), .B1(
        n8265), .Y(n1990) );
  AOI2BB2XL U9939 ( .B0(n9112), .B1(n8217), .A0N(\xArray[15][35] ), .A1N(n8256), .Y(n1119) );
  AOI2BB2XL U9940 ( .B0(n9104), .B1(n8217), .A0N(\xArray[15][36] ), .A1N(n8256), .Y(n1114) );
  OA22XL U9941 ( .A0(\xArray[14][37] ), .A1(n8272), .B0(\xArray[2][37] ), .B1(
        n8185), .Y(n1403) );
  AOI22XL U9942 ( .A0(n8060), .A1(n7399), .B0(\xArray[8][12] ), .B1(n3154), 
        .Y(n3205) );
  AOI22XL U9943 ( .A0(n8137), .A1(n7399), .B0(\xArray[2][12] ), .B1(n8134), 
        .Y(n2702) );
  AOI22XL U9944 ( .A0(n8060), .A1(n7397), .B0(\xArray[8][11] ), .B1(n8057), 
        .Y(n3206) );
  AOI22XL U9945 ( .A0(n8137), .A1(n7397), .B0(\xArray[2][11] ), .B1(n8134), 
        .Y(n2704) );
  AOI22XL U9946 ( .A0(n8060), .A1(n7395), .B0(\xArray[8][10] ), .B1(n8056), 
        .Y(n3207) );
  AOI22XL U9947 ( .A0(n8137), .A1(n7395), .B0(\xArray[2][10] ), .B1(n8134), 
        .Y(n2706) );
  OAI22XL U9948 ( .A0(\xArray[10][12] ), .A1(n7893), .B0(n7896), .B1(n7399), 
        .Y(n3348) );
  OAI22XL U9949 ( .A0(\xArray[13][12] ), .A1(n7868), .B0(n7880), .B1(n7399), 
        .Y(n3553) );
  OAI22XL U9950 ( .A0(\xArray[10][11] ), .A1(n7893), .B0(n7896), .B1(n7397), 
        .Y(n3349) );
  OAI22XL U9951 ( .A0(\xArray[13][11] ), .A1(n7868), .B0(n7884), .B1(n7397), 
        .Y(n3554) );
  OAI22XL U9952 ( .A0(\xArray[1][12] ), .A1(n7788), .B0(n7801), .B1(n7399), 
        .Y(n2581) );
  OAI22XL U9953 ( .A0(\xArray[1][11] ), .A1(n7788), .B0(n7801), .B1(n7397), 
        .Y(n2582) );
  OAI22XL U9954 ( .A0(\xArray[1][10] ), .A1(n7787), .B0(n7802), .B1(n7395), 
        .Y(n2583) );
  OAI22XL U9955 ( .A0(\xArray[10][10] ), .A1(n7893), .B0(n7895), .B1(n7395), 
        .Y(n3350) );
  OAI22XL U9956 ( .A0(\xArray[13][10] ), .A1(n7868), .B0(n7884), .B1(n7395), 
        .Y(n3555) );
  OAI22XL U9957 ( .A0(\xArray[0][12] ), .A1(n7768), .B0(n7777), .B1(n7399), 
        .Y(n2485) );
  OAI22XL U9958 ( .A0(\xArray[0][11] ), .A1(n7768), .B0(n7777), .B1(n7397), 
        .Y(n2488) );
  OAI22XL U9959 ( .A0(\xArray[0][10] ), .A1(n7768), .B0(n7777), .B1(n7395), 
        .Y(n2491) );
  OAI22XL U9960 ( .A0(\xArray[11][11] ), .A1(n7831), .B0(n7836), .B1(n7397), 
        .Y(n3417) );
  OAI22XL U9961 ( .A0(\xArray[11][10] ), .A1(n7831), .B0(n7835), .B1(n7395), 
        .Y(n3418) );
  OAI22XL U9962 ( .A0(\xArray[6][11] ), .A1(n7811), .B0(n7816), .B1(n7397), 
        .Y(n3065) );
  OAI22XL U9963 ( .A0(\xArray[6][10] ), .A1(n7811), .B0(n7815), .B1(n7395), 
        .Y(n3066) );
  OAI22XL U9964 ( .A0(\xArray[7][11] ), .A1(n7850), .B0(n7855), .B1(n7397), 
        .Y(n3136) );
  OAI22XL U9965 ( .A0(\xArray[12][11] ), .A1(n7913), .B0(n7926), .B1(n7397), 
        .Y(n3486) );
  OAI22XL U9966 ( .A0(\xArray[7][10] ), .A1(n7850), .B0(n7854), .B1(n7395), 
        .Y(n3137) );
  OAI22XL U9967 ( .A0(\xArray[12][10] ), .A1(n7913), .B0(n7918), .B1(n7395), 
        .Y(n3487) );
  OA22XL U9968 ( .A0(n8312), .A1(n1430), .B0(n7729), .B1(n1652), .Y(n2045) );
  OA22XL U9969 ( .A0(n8312), .A1(n1434), .B0(n7729), .B1(n1655), .Y(n2054) );
  MX4XL U9970 ( .A(\bArray[4][33] ), .B(\bArray[5][33] ), .C(\bArray[6][33] ), 
        .D(\bArray[7][33] ), .S0(n7210), .S1(n8409), .Y(n7078) );
  MX4XL U9971 ( .A(\bArray[12][33] ), .B(\bArray[13][33] ), .C(
        \bArray[14][33] ), .D(\bArray[15][33] ), .S0(n7210), .S1(n8409), .Y(
        n7076) );
  MX4XL U9972 ( .A(\bArray[8][33] ), .B(\bArray[9][33] ), .C(\bArray[10][33] ), 
        .D(\bArray[11][33] ), .S0(n7210), .S1(n8409), .Y(n7077) );
  MX4XL U9973 ( .A(\bArray[4][34] ), .B(\bArray[5][34] ), .C(\bArray[6][34] ), 
        .D(\bArray[7][34] ), .S0(n7200), .S1(n7222), .Y(n7082) );
  MX4XL U9974 ( .A(\bArray[12][34] ), .B(\bArray[13][34] ), .C(
        \bArray[14][34] ), .D(\bArray[15][34] ), .S0(n7200), .S1(n7222), .Y(
        n7080) );
  MX4XL U9975 ( .A(\bArray[8][34] ), .B(\bArray[9][34] ), .C(\bArray[10][34] ), 
        .D(\bArray[11][34] ), .S0(n7200), .S1(n7222), .Y(n7081) );
  INVXL U9976 ( .A(\xArray[5][23] ), .Y(n9210) );
  INVXL U9977 ( .A(\xArray[5][24] ), .Y(n9202) );
  INVXL U9978 ( .A(\xArray[14][32] ), .Y(n9142) );
  INVX1 U9979 ( .A(\xArray[14][33] ), .Y(n9134) );
  INVXL U9980 ( .A(\xArray[9][23] ), .Y(n9212) );
  INVXL U9981 ( .A(\xArray[9][24] ), .Y(n9204) );
  AOI2BB2XL U9982 ( .B0(n9110), .B1(n8203), .A0N(\xArray[10][36] ), .A1N(n8255), .Y(n1996) );
  INVXL U9983 ( .A(\xArray[3][32] ), .Y(n9136) );
  INVXL U9984 ( .A(\xArray[6][23] ), .Y(n9211) );
  INVXL U9985 ( .A(\xArray[10][23] ), .Y(n9213) );
  MX4XL U9986 ( .A(\bArray[0][33] ), .B(\bArray[1][33] ), .C(\bArray[2][33] ), 
        .D(\bArray[3][33] ), .S0(n7200), .S1(n7222), .Y(n7079) );
  OA22XL U9987 ( .A0(\xArray[14][38] ), .A1(n8270), .B0(\xArray[2][38] ), .B1(
        n8185), .Y(n1399) );
  OA22XL U9988 ( .A0(\xArray[15][38] ), .A1(n8193), .B0(\xArray[11][38] ), 
        .B1(n8264), .Y(n1980) );
  OA22XL U9989 ( .A0(\xArray[15][37] ), .A1(n8193), .B0(\xArray[11][37] ), 
        .B1(n8264), .Y(n1989) );
  OA22XL U9990 ( .A0(\xArray[4][35] ), .A1(n8197), .B0(\xArray[0][35] ), .B1(
        n8263), .Y(n1118) );
  OA22XL U9991 ( .A0(\xArray[4][36] ), .A1(n8197), .B0(\xArray[0][36] ), .B1(
        n8263), .Y(n1113) );
  OA22XL U9992 ( .A0(\xArray[5][35] ), .A1(n8195), .B0(\xArray[1][35] ), .B1(
        n8267), .Y(n870) );
  OA22XL U9993 ( .A0(\xArray[5][34] ), .A1(n8195), .B0(\xArray[1][34] ), .B1(
        n8267), .Y(n873) );
  AOI2BB2XL U9994 ( .B0(n9094), .B1(n8203), .A0N(\xArray[10][38] ), .A1N(n8254), .Y(n1978) );
  AOI2BB2XL U9995 ( .B0(n9086), .B1(n8207), .A0N(\xArray[10][39] ), .A1N(n8254), .Y(n1969) );
  AOI2BB2XL U9996 ( .B0(n9096), .B1(n8208), .A0N(\xArray[15][37] ), .A1N(n8256), .Y(n1109) );
  AOI22XL U9997 ( .A0(n8060), .A1(n7393), .B0(\xArray[8][9] ), .B1(n3154), .Y(
        n3208) );
  AOI22XL U9998 ( .A0(n8137), .A1(n7393), .B0(\xArray[2][9] ), .B1(n8134), .Y(
        n2708) );
  AOI22XL U9999 ( .A0(n8060), .A1(n7391), .B0(\xArray[8][8] ), .B1(n3154), .Y(
        n3209) );
  AOI22XL U10000 ( .A0(n8137), .A1(n7391), .B0(\xArray[2][8] ), .B1(n8134), 
        .Y(n2710) );
  AOI22XL U10001 ( .A0(n8060), .A1(n7389), .B0(\xArray[8][7] ), .B1(n3154), 
        .Y(n3210) );
  AOI22XL U10002 ( .A0(n8137), .A1(n7389), .B0(\xArray[2][7] ), .B1(n8134), 
        .Y(n2712) );
  OAI22XL U10003 ( .A0(\xArray[1][9] ), .A1(n7787), .B0(n7801), .B1(n7393), 
        .Y(n2584) );
  OAI22XL U10004 ( .A0(\xArray[10][9] ), .A1(n7893), .B0(n7895), .B1(n7393), 
        .Y(n3351) );
  OAI22XL U10005 ( .A0(\xArray[13][9] ), .A1(n7868), .B0(n7884), .B1(n7393), 
        .Y(n3556) );
  OAI22XL U10006 ( .A0(\xArray[1][8] ), .A1(n7786), .B0(n7801), .B1(n7391), 
        .Y(n2585) );
  OAI22XL U10007 ( .A0(\xArray[10][8] ), .A1(n7893), .B0(n7895), .B1(n7391), 
        .Y(n3352) );
  OAI22XL U10008 ( .A0(\xArray[13][8] ), .A1(n7868), .B0(n7884), .B1(n7391), 
        .Y(n3557) );
  OAI22XL U10009 ( .A0(\xArray[1][7] ), .A1(n7787), .B0(n7801), .B1(n7389), 
        .Y(n2586) );
  OAI22XL U10010 ( .A0(\xArray[10][7] ), .A1(n7893), .B0(n7895), .B1(n7389), 
        .Y(n3353) );
  OAI22XL U10011 ( .A0(\xArray[13][7] ), .A1(n7868), .B0(n7885), .B1(n7389), 
        .Y(n3558) );
  OAI22XL U10012 ( .A0(\xArray[0][9] ), .A1(n7768), .B0(n7778), .B1(n7393), 
        .Y(n2494) );
  OAI22XL U10013 ( .A0(\xArray[0][8] ), .A1(n7768), .B0(n7778), .B1(n7391), 
        .Y(n2497) );
  OAI22XL U10014 ( .A0(\xArray[0][7] ), .A1(n7768), .B0(n7778), .B1(n7389), 
        .Y(n2500) );
  OAI22XL U10015 ( .A0(\xArray[11][9] ), .A1(n7831), .B0(n7835), .B1(n7393), 
        .Y(n3419) );
  OAI22XL U10016 ( .A0(\xArray[11][8] ), .A1(n7831), .B0(n7835), .B1(n7391), 
        .Y(n3420) );
  OAI22XL U10017 ( .A0(\xArray[11][7] ), .A1(n7831), .B0(n7835), .B1(n7389), 
        .Y(n3421) );
  OAI22XL U10018 ( .A0(\xArray[6][9] ), .A1(n7811), .B0(n7815), .B1(n7393), 
        .Y(n3067) );
  OAI22XL U10019 ( .A0(\xArray[6][8] ), .A1(n7811), .B0(n7815), .B1(n7391), 
        .Y(n3068) );
  OAI22XL U10020 ( .A0(\xArray[6][7] ), .A1(n7811), .B0(n7815), .B1(n7389), 
        .Y(n3069) );
  OAI22XL U10021 ( .A0(\xArray[7][9] ), .A1(n7850), .B0(n7854), .B1(n7393), 
        .Y(n3138) );
  OAI22XL U10022 ( .A0(\xArray[12][9] ), .A1(n7913), .B0(n7916), .B1(n7393), 
        .Y(n3488) );
  OAI22XL U10023 ( .A0(\xArray[7][8] ), .A1(n7850), .B0(n7854), .B1(n7391), 
        .Y(n3139) );
  OAI22XL U10024 ( .A0(\xArray[12][8] ), .A1(n7913), .B0(n7916), .B1(n7391), 
        .Y(n3489) );
  OAI22XL U10025 ( .A0(\xArray[7][7] ), .A1(n7850), .B0(n7854), .B1(n7389), 
        .Y(n3140) );
  OAI22XL U10026 ( .A0(\xArray[12][7] ), .A1(n7913), .B0(n7918), .B1(n7389), 
        .Y(n3490) );
  OA22XL U10027 ( .A0(n8312), .A1(n1426), .B0(n7730), .B1(n1649), .Y(n2036) );
  OA22XL U10028 ( .A0(n8312), .A1(n1422), .B0(n7730), .B1(n1646), .Y(n2027) );
  MX4XL U10029 ( .A(\bArray[4][35] ), .B(\bArray[5][35] ), .C(\bArray[6][35] ), 
        .D(\bArray[7][35] ), .S0(n7204), .S1(N1762), .Y(n7086) );
  MX4XL U10030 ( .A(\bArray[12][35] ), .B(\bArray[13][35] ), .C(
        \bArray[14][35] ), .D(\bArray[15][35] ), .S0(n7205), .S1(n7213), .Y(
        n7084) );
  MX4XL U10031 ( .A(\bArray[8][35] ), .B(\bArray[9][35] ), .C(\bArray[10][35] ), .D(\bArray[11][35] ), .S0(n7204), .S1(N1762), .Y(n7085) );
  MX4XL U10032 ( .A(\bArray[4][36] ), .B(\bArray[5][36] ), .C(\bArray[6][36] ), 
        .D(\bArray[7][36] ), .S0(n7204), .S1(N1762), .Y(n7090) );
  MX4XL U10033 ( .A(\bArray[12][36] ), .B(\bArray[13][36] ), .C(
        \bArray[14][36] ), .D(\bArray[15][36] ), .S0(n7204), .S1(N1762), .Y(
        n7088) );
  MX4XL U10034 ( .A(\bArray[8][36] ), .B(\bArray[9][36] ), .C(\bArray[10][36] ), .D(\bArray[11][36] ), .S0(n7204), .S1(N1762), .Y(n7089) );
  INVXL U10035 ( .A(\xArray[5][25] ), .Y(n9194) );
  INVXL U10036 ( .A(\xArray[5][26] ), .Y(n9186) );
  INVX1 U10037 ( .A(\xArray[14][34] ), .Y(n9126) );
  INVX1 U10038 ( .A(\xArray[14][35] ), .Y(n9118) );
  INVXL U10039 ( .A(\xArray[9][25] ), .Y(n9196) );
  INVXL U10040 ( .A(\xArray[9][26] ), .Y(n9188) );
  INVXL U10041 ( .A(\xArray[3][33] ), .Y(n9128) );
  INVXL U10042 ( .A(\xArray[3][34] ), .Y(n9120) );
  INVXL U10043 ( .A(\xArray[6][24] ), .Y(n9203) );
  INVXL U10044 ( .A(\xArray[6][25] ), .Y(n9195) );
  INVXL U10045 ( .A(\xArray[10][24] ), .Y(n9205) );
  INVXL U10046 ( .A(\xArray[10][25] ), .Y(n9197) );
  MX4XL U10047 ( .A(\bArray[0][35] ), .B(\bArray[1][35] ), .C(\bArray[2][35] ), 
        .D(\bArray[3][35] ), .S0(n7204), .S1(N1762), .Y(n7087) );
  MX4XL U10048 ( .A(\bArray[0][36] ), .B(\bArray[1][36] ), .C(\bArray[2][36] ), 
        .D(\bArray[3][36] ), .S0(n7204), .S1(N1762), .Y(n7091) );
  OA22XL U10049 ( .A0(\xArray[14][39] ), .A1(n8271), .B0(\xArray[2][39] ), 
        .B1(n8185), .Y(n1395) );
  OA22XL U10050 ( .A0(\xArray[14][40] ), .A1(n8270), .B0(\xArray[2][40] ), 
        .B1(n8185), .Y(n1391) );
  OA22XL U10051 ( .A0(\xArray[0][39] ), .A1(n8193), .B0(\xArray[12][39] ), 
        .B1(n8264), .Y(n1972) );
  OA22XL U10052 ( .A0(\xArray[15][39] ), .A1(n8193), .B0(\xArray[11][39] ), 
        .B1(n8264), .Y(n1971) );
  OA22XL U10053 ( .A0(\xArray[4][37] ), .A1(n8197), .B0(\xArray[0][37] ), .B1(
        n8263), .Y(n1108) );
  OA22XL U10054 ( .A0(\xArray[0][40] ), .A1(n8193), .B0(\xArray[12][40] ), 
        .B1(n8264), .Y(n1963) );
  OA22XL U10055 ( .A0(\xArray[15][40] ), .A1(n8193), .B0(\xArray[11][40] ), 
        .B1(n8264), .Y(n1962) );
  OA22XL U10056 ( .A0(\xArray[5][36] ), .A1(n8195), .B0(\xArray[1][36] ), .B1(
        n8267), .Y(n867) );
  OA22XL U10057 ( .A0(\xArray[5][39] ), .A1(n8194), .B0(\xArray[1][39] ), .B1(
        n8265), .Y(n858) );
  AOI2BB2XL U10058 ( .B0(n9078), .B1(n8212), .A0N(\xArray[10][40] ), .A1N(
        n8254), .Y(n1960) );
  OA22XL U10059 ( .A0(\xArray[14][41] ), .A1(n8271), .B0(\xArray[2][41] ), 
        .B1(n8185), .Y(n1387) );
  AOI22XL U10060 ( .A0(n8060), .A1(n7387), .B0(\xArray[8][6] ), .B1(n3154), 
        .Y(n3211) );
  AOI22XL U10061 ( .A0(n8137), .A1(n7387), .B0(\xArray[2][6] ), .B1(n8134), 
        .Y(n2714) );
  AOI22XL U10062 ( .A0(n8060), .A1(n7385), .B0(\xArray[8][5] ), .B1(n3154), 
        .Y(n3212) );
  AOI22XL U10063 ( .A0(n8137), .A1(n7385), .B0(\xArray[2][5] ), .B1(n8134), 
        .Y(n2716) );
  AOI22XL U10064 ( .A0(n8060), .A1(n7383), .B0(\xArray[8][4] ), .B1(n3154), 
        .Y(n3213) );
  AOI22XL U10065 ( .A0(n8137), .A1(n7383), .B0(\xArray[2][4] ), .B1(n8134), 
        .Y(n2718) );
  OAI22XL U10066 ( .A0(\xArray[1][6] ), .A1(n7786), .B0(n7802), .B1(n7387), 
        .Y(n2587) );
  OAI22XL U10067 ( .A0(\xArray[10][6] ), .A1(n7893), .B0(n7897), .B1(n7387), 
        .Y(n3354) );
  OAI22XL U10068 ( .A0(\xArray[13][6] ), .A1(n7868), .B0(n7885), .B1(n7387), 
        .Y(n3559) );
  OAI22XL U10069 ( .A0(\xArray[1][5] ), .A1(n7786), .B0(n7802), .B1(n7385), 
        .Y(n2588) );
  OAI22XL U10070 ( .A0(\xArray[10][5] ), .A1(n7893), .B0(n7900), .B1(n7385), 
        .Y(n3355) );
  OAI22XL U10071 ( .A0(\xArray[13][5] ), .A1(n7868), .B0(n7885), .B1(n7385), 
        .Y(n3560) );
  OAI22XL U10072 ( .A0(\xArray[1][4] ), .A1(n7786), .B0(n7802), .B1(n7383), 
        .Y(n2589) );
  OAI22XL U10073 ( .A0(\xArray[10][4] ), .A1(n7893), .B0(n7897), .B1(n7383), 
        .Y(n3356) );
  OAI22XL U10074 ( .A0(\xArray[13][4] ), .A1(n7868), .B0(n7885), .B1(n7383), 
        .Y(n3561) );
  OAI22XL U10075 ( .A0(\xArray[0][6] ), .A1(n7768), .B0(n7778), .B1(n7387), 
        .Y(n2503) );
  OAI22XL U10076 ( .A0(\xArray[0][5] ), .A1(n7768), .B0(n7777), .B1(n7385), 
        .Y(n2506) );
  OAI22XL U10077 ( .A0(\xArray[0][4] ), .A1(n7768), .B0(n7777), .B1(n7383), 
        .Y(n2509) );
  OAI22XL U10078 ( .A0(\xArray[11][6] ), .A1(n7831), .B0(n7844), .B1(n7387), 
        .Y(n3422) );
  OAI22XL U10079 ( .A0(\xArray[11][5] ), .A1(n7831), .B0(n7836), .B1(n7385), 
        .Y(n3423) );
  OAI22XL U10080 ( .A0(\xArray[11][4] ), .A1(n7831), .B0(n7836), .B1(n7383), 
        .Y(n3424) );
  OAI22XL U10081 ( .A0(\xArray[6][6] ), .A1(n7811), .B0(n7814), .B1(n7387), 
        .Y(n3070) );
  OAI22XL U10082 ( .A0(\xArray[6][5] ), .A1(n7811), .B0(n7816), .B1(n7385), 
        .Y(n3071) );
  OAI22XL U10083 ( .A0(\xArray[6][4] ), .A1(n7811), .B0(n7816), .B1(n7383), 
        .Y(n3072) );
  OAI22XL U10084 ( .A0(\xArray[7][6] ), .A1(n7850), .B0(n7855), .B1(n7387), 
        .Y(n3141) );
  OAI22XL U10085 ( .A0(\xArray[12][6] ), .A1(n7913), .B0(n7916), .B1(n7387), 
        .Y(n3491) );
  OAI22XL U10086 ( .A0(\xArray[7][5] ), .A1(n7850), .B0(n7855), .B1(n7385), 
        .Y(n3142) );
  OAI22XL U10087 ( .A0(\xArray[12][5] ), .A1(n7913), .B0(n7915), .B1(n7385), 
        .Y(n3492) );
  OAI22XL U10088 ( .A0(\xArray[7][4] ), .A1(n7850), .B0(n7855), .B1(n7383), 
        .Y(n3143) );
  OAI22XL U10089 ( .A0(\xArray[12][4] ), .A1(n7913), .B0(n7916), .B1(n7383), 
        .Y(n3493) );
  OA22XL U10090 ( .A0(n8312), .A1(n1418), .B0(n7730), .B1(n1643), .Y(n2018) );
  OA22XL U10091 ( .A0(n8312), .A1(n1414), .B0(n7730), .B1(n1640), .Y(n2009) );
  MX4XL U10092 ( .A(\bArray[4][37] ), .B(\bArray[5][37] ), .C(\bArray[6][37] ), 
        .D(\bArray[7][37] ), .S0(n7204), .S1(N1762), .Y(n7094) );
  MX4XL U10093 ( .A(\bArray[12][37] ), .B(\bArray[13][37] ), .C(
        \bArray[14][37] ), .D(\bArray[15][37] ), .S0(n7204), .S1(N1762), .Y(
        n7092) );
  MX4XL U10094 ( .A(\bArray[8][37] ), .B(\bArray[9][37] ), .C(\bArray[10][37] ), .D(\bArray[11][37] ), .S0(n7204), .S1(N1762), .Y(n7093) );
  INVXL U10095 ( .A(\xArray[5][27] ), .Y(n9178) );
  INVXL U10096 ( .A(\xArray[5][28] ), .Y(n9170) );
  AOI2BB2XL U10097 ( .B0(n9080), .B1(n8214), .A0N(\xArray[15][39] ), .A1N(
        n8256), .Y(n1099) );
  AOI2BB2XL U10098 ( .B0(n9072), .B1(n8208), .A0N(\xArray[15][40] ), .A1N(
        n8256), .Y(n1094) );
  INVX1 U10099 ( .A(\xArray[14][36] ), .Y(n9110) );
  INVX1 U10100 ( .A(\xArray[14][37] ), .Y(n9102) );
  INVXL U10101 ( .A(\xArray[9][27] ), .Y(n9180) );
  INVXL U10102 ( .A(\xArray[9][28] ), .Y(n9172) );
  INVXL U10103 ( .A(\xArray[3][35] ), .Y(n9112) );
  INVXL U10104 ( .A(\xArray[3][36] ), .Y(n9104) );
  INVXL U10105 ( .A(\xArray[6][26] ), .Y(n9187) );
  INVXL U10106 ( .A(\xArray[6][27] ), .Y(n9179) );
  INVXL U10107 ( .A(\xArray[10][26] ), .Y(n9189) );
  INVXL U10108 ( .A(\xArray[10][27] ), .Y(n9181) );
  MX4XL U10109 ( .A(\bArray[0][37] ), .B(\bArray[1][37] ), .C(\bArray[2][37] ), 
        .D(\bArray[3][37] ), .S0(n7204), .S1(N1762), .Y(n7095) );
  OA22XL U10110 ( .A0(\xArray[4][39] ), .A1(n8183), .B0(\xArray[0][39] ), .B1(
        n8254), .Y(n1098) );
  OA22XL U10111 ( .A0(\xArray[0][41] ), .A1(n8193), .B0(\xArray[12][41] ), 
        .B1(n8264), .Y(n1954) );
  OA22XL U10112 ( .A0(\xArray[15][41] ), .A1(n8193), .B0(\xArray[11][41] ), 
        .B1(n8264), .Y(n1953) );
  OA22XL U10113 ( .A0(\xArray[4][40] ), .A1(n8183), .B0(\xArray[0][40] ), .B1(
        n8254), .Y(n1093) );
  OA22XL U10114 ( .A0(\xArray[0][42] ), .A1(n8193), .B0(\xArray[12][42] ), 
        .B1(n8263), .Y(n1945) );
  OA22XL U10115 ( .A0(\xArray[15][42] ), .A1(n8193), .B0(\xArray[11][42] ), 
        .B1(n8267), .Y(n1944) );
  AOI2BB2XL U10116 ( .B0(n9062), .B1(n8203), .A0N(\xArray[10][42] ), .A1N(
        n8254), .Y(n1942) );
  AOI2BB2XL U10117 ( .B0(n9070), .B1(n8208), .A0N(\xArray[10][41] ), .A1N(
        n8254), .Y(n1951) );
  AOI2BB2XL U10118 ( .B0(n9064), .B1(n8214), .A0N(\xArray[15][41] ), .A1N(
        n8257), .Y(n1089) );
  OA22XL U10119 ( .A0(\xArray[1][43] ), .A1(n8199), .B0(\xArray[13][43] ), 
        .B1(n8269), .Y(n1614) );
  AOI22XL U10120 ( .A0(n8060), .A1(n7381), .B0(\xArray[8][3] ), .B1(n8056), 
        .Y(n3214) );
  AOI22XL U10121 ( .A0(n8137), .A1(n7381), .B0(\xArray[2][3] ), .B1(n8133), 
        .Y(n2720) );
  AOI22XL U10122 ( .A0(n8060), .A1(n7379), .B0(\xArray[8][2] ), .B1(n8056), 
        .Y(n3215) );
  AOI22XL U10123 ( .A0(n8137), .A1(n7379), .B0(\xArray[2][2] ), .B1(n8132), 
        .Y(n2722) );
  AOI22XL U10124 ( .A0(n8060), .A1(n7377), .B0(\xArray[8][1] ), .B1(n8055), 
        .Y(n3216) );
  AOI22XL U10125 ( .A0(n8137), .A1(n7377), .B0(\xArray[2][1] ), .B1(n8133), 
        .Y(n2724) );
  OAI22XL U10126 ( .A0(\xArray[1][3] ), .A1(n7785), .B0(n7802), .B1(n7381), 
        .Y(n2590) );
  OAI22XL U10127 ( .A0(\xArray[10][3] ), .A1(n7894), .B0(n7908), .B1(n7381), 
        .Y(n3357) );
  OAI22XL U10128 ( .A0(\xArray[13][3] ), .A1(n7868), .B0(n7884), .B1(n7381), 
        .Y(n3562) );
  OAI22XL U10129 ( .A0(\xArray[1][2] ), .A1(n7785), .B0(n7803), .B1(n7379), 
        .Y(n2591) );
  OAI22XL U10130 ( .A0(\xArray[10][2] ), .A1(n7894), .B0(n7897), .B1(n7379), 
        .Y(n3358) );
  OAI22XL U10131 ( .A0(\xArray[13][2] ), .A1(n7868), .B0(n7885), .B1(n7379), 
        .Y(n3563) );
  OAI22XL U10132 ( .A0(\xArray[1][1] ), .A1(n7785), .B0(n7803), .B1(n7377), 
        .Y(n2592) );
  OAI22XL U10133 ( .A0(\xArray[10][1] ), .A1(n7894), .B0(n7908), .B1(n7377), 
        .Y(n3359) );
  OAI22XL U10134 ( .A0(\xArray[13][1] ), .A1(n7868), .B0(n7885), .B1(n7377), 
        .Y(n3564) );
  OAI22XL U10135 ( .A0(\xArray[0][3] ), .A1(n7768), .B0(n7777), .B1(n7381), 
        .Y(n2512) );
  OAI22XL U10136 ( .A0(\xArray[0][2] ), .A1(n7768), .B0(n7778), .B1(n7379), 
        .Y(n2515) );
  OAI22XL U10137 ( .A0(\xArray[0][1] ), .A1(n7768), .B0(n7778), .B1(n7377), 
        .Y(n2518) );
  OAI22XL U10138 ( .A0(\xArray[11][3] ), .A1(n7832), .B0(n7834), .B1(n7381), 
        .Y(n3425) );
  OAI22XL U10139 ( .A0(\xArray[11][2] ), .A1(n7832), .B0(n7833), .B1(n7379), 
        .Y(n3426) );
  OAI22XL U10140 ( .A0(\xArray[11][1] ), .A1(n7832), .B0(n7844), .B1(n7377), 
        .Y(n3427) );
  OAI22XL U10141 ( .A0(\xArray[6][3] ), .A1(n7812), .B0(n7816), .B1(n7381), 
        .Y(n3073) );
  OAI22XL U10142 ( .A0(\xArray[6][2] ), .A1(n7812), .B0(n7813), .B1(n7379), 
        .Y(n3074) );
  OAI22XL U10143 ( .A0(\xArray[6][1] ), .A1(n7812), .B0(n7823), .B1(n7377), 
        .Y(n3075) );
  OAI22XL U10144 ( .A0(\xArray[7][3] ), .A1(n7851), .B0(n7853), .B1(n7381), 
        .Y(n3144) );
  OAI22XL U10145 ( .A0(\xArray[12][3] ), .A1(n7914), .B0(n7915), .B1(n7381), 
        .Y(n3494) );
  OAI22XL U10146 ( .A0(\xArray[7][2] ), .A1(n7851), .B0(n7852), .B1(n7379), 
        .Y(n3145) );
  OAI22XL U10147 ( .A0(\xArray[12][2] ), .A1(n7914), .B0(n7916), .B1(n7379), 
        .Y(n3495) );
  OAI22XL U10148 ( .A0(\xArray[7][1] ), .A1(n7851), .B0(n7857), .B1(n7377), 
        .Y(n3146) );
  OAI22XL U10149 ( .A0(\xArray[12][1] ), .A1(n7914), .B0(n7926), .B1(n7377), 
        .Y(n3496) );
  OA22XL U10150 ( .A0(n8312), .A1(n1410), .B0(n7730), .B1(n1637), .Y(n2000) );
  OA22XL U10151 ( .A0(n8310), .A1(n1406), .B0(n7730), .B1(n1634), .Y(n1991) );
  MX4XL U10152 ( .A(\bArray[4][39] ), .B(\bArray[5][39] ), .C(\bArray[6][39] ), 
        .D(\bArray[7][39] ), .S0(n7209), .S1(n7219), .Y(n7102) );
  MX4XL U10153 ( .A(\bArray[12][39] ), .B(\bArray[13][39] ), .C(
        \bArray[14][39] ), .D(\bArray[15][39] ), .S0(n7205), .S1(N1762), .Y(
        n7100) );
  MX4XL U10154 ( .A(\bArray[8][39] ), .B(\bArray[9][39] ), .C(\bArray[10][39] ), .D(\bArray[11][39] ), .S0(n7200), .S1(n7222), .Y(n7101) );
  MX4XL U10155 ( .A(\bArray[4][40] ), .B(\bArray[5][40] ), .C(\bArray[6][40] ), 
        .D(\bArray[7][40] ), .S0(n7200), .S1(n7215), .Y(n7106) );
  MX4XL U10156 ( .A(\bArray[12][40] ), .B(\bArray[13][40] ), .C(
        \bArray[14][40] ), .D(\bArray[15][40] ), .S0(n7206), .S1(n7219), .Y(
        n7104) );
  MX4XL U10157 ( .A(\bArray[8][40] ), .B(\bArray[9][40] ), .C(\bArray[10][40] ), .D(\bArray[11][40] ), .S0(n7205), .S1(n7219), .Y(n7105) );
  INVXL U10158 ( .A(\xArray[5][29] ), .Y(n9162) );
  INVXL U10159 ( .A(\xArray[5][30] ), .Y(n9154) );
  INVXL U10160 ( .A(\xArray[9][29] ), .Y(n9164) );
  INVXL U10161 ( .A(\xArray[9][30] ), .Y(n9156) );
  INVXL U10162 ( .A(\xArray[3][37] ), .Y(n9096) );
  INVXL U10163 ( .A(\xArray[3][38] ), .Y(n9088) );
  INVXL U10164 ( .A(\xArray[6][28] ), .Y(n9171) );
  INVXL U10165 ( .A(\xArray[6][29] ), .Y(n9163) );
  INVXL U10166 ( .A(\xArray[10][28] ), .Y(n9173) );
  INVXL U10167 ( .A(\xArray[10][29] ), .Y(n9165) );
  MX4XL U10168 ( .A(\bArray[0][39] ), .B(\bArray[1][39] ), .C(\bArray[2][39] ), 
        .D(\bArray[3][39] ), .S0(n7207), .S1(n7219), .Y(n7103) );
  MX4XL U10169 ( .A(\bArray[0][40] ), .B(\bArray[1][40] ), .C(\bArray[2][40] ), 
        .D(\bArray[3][40] ), .S0(n7210), .S1(n7215), .Y(n7107) );
  OA22XL U10170 ( .A0(\xArray[1][42] ), .A1(n8199), .B0(\xArray[13][42] ), 
        .B1(n8254), .Y(n1617) );
  OA22XL U10171 ( .A0(\xArray[4][41] ), .A1(n8183), .B0(\xArray[0][41] ), .B1(
        n8254), .Y(n1088) );
  OA22XL U10172 ( .A0(\xArray[0][43] ), .A1(n8193), .B0(\xArray[12][43] ), 
        .B1(n8263), .Y(n1936) );
  OA22XL U10173 ( .A0(\xArray[15][43] ), .A1(n8193), .B0(\xArray[11][43] ), 
        .B1(n8263), .Y(n1935) );
  OA22XL U10174 ( .A0(\xArray[14][42] ), .A1(n8270), .B0(\xArray[2][42] ), 
        .B1(n8185), .Y(n1383) );
  OA22XL U10175 ( .A0(\xArray[4][42] ), .A1(n6707), .B0(\xArray[0][42] ), .B1(
        n8254), .Y(n1083) );
  OA22XL U10176 ( .A0(\xArray[0][44] ), .A1(n8193), .B0(\xArray[12][44] ), 
        .B1(n8263), .Y(n1927) );
  OA22XL U10177 ( .A0(\xArray[15][44] ), .A1(n8193), .B0(\xArray[11][44] ), 
        .B1(n8263), .Y(n1926) );
  OA22XL U10178 ( .A0(\xArray[14][43] ), .A1(n8271), .B0(\xArray[2][43] ), 
        .B1(n8185), .Y(n1379) );
  OA22XL U10179 ( .A0(\xArray[5][40] ), .A1(n8194), .B0(\xArray[1][40] ), .B1(
        n8271), .Y(n855) );
  OA22XL U10180 ( .A0(\xArray[5][41] ), .A1(n8194), .B0(\xArray[1][41] ), .B1(
        n8255), .Y(n852) );
  AOI2BB2XL U10181 ( .B0(n9054), .B1(n8217), .A0N(\xArray[10][43] ), .A1N(
        n8254), .Y(n1933) );
  AOI2BB2XL U10182 ( .B0(n9046), .B1(n8217), .A0N(\xArray[10][44] ), .A1N(
        n8254), .Y(n1924) );
  AOI2BB2XL U10183 ( .B0(n9038), .B1(n8217), .A0N(\xArray[10][45] ), .A1N(
        n8254), .Y(n1915) );
  AOI2BB2XL U10184 ( .B0(n9030), .B1(n8216), .A0N(\xArray[10][46] ), .A1N(
        n8254), .Y(n1906) );
  OA22XL U10185 ( .A0(\xArray[0][47] ), .A1(n8199), .B0(\xArray[12][47] ), 
        .B1(n8263), .Y(n1900) );
  AOI2BB2XL U10186 ( .B0(n9056), .B1(n8208), .A0N(\xArray[15][42] ), .A1N(
        n8257), .Y(n1084) );
  AOI2BB2XL U10187 ( .B0(n9048), .B1(n8217), .A0N(\xArray[15][43] ), .A1N(
        n8257), .Y(n1079) );
  AOI2BB2XL U10188 ( .B0(n9040), .B1(n8217), .A0N(\xArray[15][44] ), .A1N(
        n8257), .Y(n1074) );
  OA22XL U10189 ( .A0(\xArray[14][47] ), .A1(n8272), .B0(\xArray[2][47] ), 
        .B1(n8184), .Y(n1363) );
  OA22XL U10190 ( .A0(\xArray[4][45] ), .A1(n8196), .B0(\xArray[0][45] ), .B1(
        n8254), .Y(n1068) );
  OA22XL U10191 ( .A0(\xArray[14][46] ), .A1(n8273), .B0(\xArray[2][46] ), 
        .B1(n8184), .Y(n1367) );
  OA22XL U10192 ( .A0(\xArray[15][46] ), .A1(n8193), .B0(\xArray[11][46] ), 
        .B1(n8263), .Y(n1908) );
  OA22XL U10193 ( .A0(\xArray[15][47] ), .A1(n8193), .B0(\xArray[11][47] ), 
        .B1(n8263), .Y(n1899) );
  OA22XL U10194 ( .A0(\xArray[1][44] ), .A1(n8199), .B0(\xArray[13][44] ), 
        .B1(n8254), .Y(n1611) );
  OA22XL U10195 ( .A0(\xArray[1][45] ), .A1(n8199), .B0(\xArray[13][45] ), 
        .B1(n8256), .Y(n1608) );
  OA22XL U10196 ( .A0(\xArray[1][46] ), .A1(n8199), .B0(\xArray[13][46] ), 
        .B1(n8256), .Y(n1605) );
  OA22XL U10197 ( .A0(\xArray[1][47] ), .A1(n8199), .B0(\xArray[13][47] ), 
        .B1(n8266), .Y(n1602) );
  AOI22XL U10198 ( .A0(n8060), .A1(n7375), .B0(\xArray[8][0] ), .B1(n8057), 
        .Y(n3217) );
  AOI22XL U10199 ( .A0(n8137), .A1(n7375), .B0(\xArray[2][0] ), .B1(n8134), 
        .Y(n2726) );
  OAI22XL U10200 ( .A0(\xArray[1][0] ), .A1(n7785), .B0(n7803), .B1(n7375), 
        .Y(n2593) );
  OAI22XL U10201 ( .A0(\xArray[10][0] ), .A1(n7894), .B0(n7900), .B1(n7375), 
        .Y(n3360) );
  OAI22XL U10202 ( .A0(\xArray[13][0] ), .A1(n7868), .B0(n7884), .B1(n7375), 
        .Y(n3565) );
  OAI22XL U10203 ( .A0(\xArray[0][0] ), .A1(n7768), .B0(n7778), .B1(n7375), 
        .Y(n2521) );
  OAI22XL U10204 ( .A0(\xArray[11][0] ), .A1(n7832), .B0(n7839), .B1(n7375), 
        .Y(n3428) );
  OAI22XL U10205 ( .A0(\xArray[6][0] ), .A1(n7812), .B0(n7819), .B1(n7375), 
        .Y(n3076) );
  OAI22XL U10206 ( .A0(\xArray[7][0] ), .A1(n7851), .B0(n7859), .B1(n7375), 
        .Y(n3147) );
  OAI22XL U10207 ( .A0(\xArray[12][0] ), .A1(n7914), .B0(n7920), .B1(n7375), 
        .Y(n3497) );
  OA22XL U10208 ( .A0(n8310), .A1(n1402), .B0(n7730), .B1(n1631), .Y(n1982) );
  OA22XL U10209 ( .A0(n8310), .A1(n1398), .B0(n7730), .B1(n1628), .Y(n1973) );
  OA22XL U10210 ( .A0(n8310), .A1(n1394), .B0(n7730), .B1(n1625), .Y(n1964) );
  MX4XL U10211 ( .A(\bArray[12][41] ), .B(\bArray[13][41] ), .C(
        \bArray[14][41] ), .D(\bArray[15][41] ), .S0(n7210), .S1(n7215), .Y(
        n7108) );
  MX4XL U10212 ( .A(\bArray[4][42] ), .B(\bArray[5][42] ), .C(\bArray[6][42] ), 
        .D(\bArray[7][42] ), .S0(n8410), .S1(n7215), .Y(n7114) );
  MX4XL U10213 ( .A(\bArray[12][42] ), .B(\bArray[13][42] ), .C(
        \bArray[14][42] ), .D(\bArray[15][42] ), .S0(n8410), .S1(n7215), .Y(
        n7112) );
  MX4XL U10214 ( .A(\bArray[8][42] ), .B(\bArray[9][42] ), .C(\bArray[10][42] ), .D(\bArray[11][42] ), .S0(n8410), .S1(n7215), .Y(n7113) );
  MX4XL U10215 ( .A(\bArray[4][43] ), .B(\bArray[5][43] ), .C(\bArray[6][43] ), 
        .D(\bArray[7][43] ), .S0(n8410), .S1(n7219), .Y(n7118) );
  MX4XL U10216 ( .A(\bArray[12][43] ), .B(\bArray[13][43] ), .C(
        \bArray[14][43] ), .D(\bArray[15][43] ), .S0(n8410), .S1(n7215), .Y(
        n7116) );
  MX4XL U10217 ( .A(\bArray[8][43] ), .B(\bArray[9][43] ), .C(\bArray[10][43] ), .D(\bArray[11][43] ), .S0(n8410), .S1(n7215), .Y(n7117) );
  INVXL U10218 ( .A(\xArray[5][31] ), .Y(n9146) );
  AOI2BB2XL U10219 ( .B0(n9032), .B1(n8217), .A0N(\xArray[15][45] ), .A1N(
        n8257), .Y(n1069) );
  INVX1 U10220 ( .A(\xArray[14][41] ), .Y(n9070) );
  INVXL U10221 ( .A(\xArray[5][32] ), .Y(n9138) );
  INVXL U10222 ( .A(\xArray[5][33] ), .Y(n9130) );
  INVXL U10223 ( .A(\xArray[5][34] ), .Y(n9122) );
  INVXL U10224 ( .A(\xArray[9][31] ), .Y(n9148) );
  INVXL U10225 ( .A(\xArray[3][39] ), .Y(n9080) );
  INVXL U10226 ( .A(\xArray[3][40] ), .Y(n9072) );
  INVXL U10227 ( .A(\xArray[3][41] ), .Y(n9064) );
  NAND2BX1 U10228 ( .AN(n456), .B(n457), .Y(N34065) );
  NAND2BX1 U10229 ( .AN(n464), .B(n465), .Y(N34064) );
  INVXL U10230 ( .A(\xArray[9][32] ), .Y(n9140) );
  INVXL U10231 ( .A(\xArray[9][33] ), .Y(n9132) );
  INVXL U10232 ( .A(\xArray[9][34] ), .Y(n9124) );
  INVXL U10233 ( .A(\xArray[6][30] ), .Y(n9155) );
  INVXL U10234 ( .A(\xArray[6][31] ), .Y(n9147) );
  INVXL U10235 ( .A(\xArray[10][30] ), .Y(n9157) );
  INVXL U10236 ( .A(\xArray[10][31] ), .Y(n9149) );
  INVXL U10237 ( .A(\xArray[6][33] ), .Y(n9131) );
  INVXL U10238 ( .A(\xArray[6][32] ), .Y(n9139) );
  INVXL U10239 ( .A(\xArray[10][33] ), .Y(n9133) );
  INVXL U10240 ( .A(\xArray[10][32] ), .Y(n9141) );
  MX4XL U10241 ( .A(\bArray[0][42] ), .B(\bArray[1][42] ), .C(\bArray[2][42] ), 
        .D(\bArray[3][42] ), .S0(n8410), .S1(n7215), .Y(n7115) );
  MX4XL U10242 ( .A(\bArray[0][43] ), .B(\bArray[1][43] ), .C(\bArray[2][43] ), 
        .D(\bArray[3][43] ), .S0(n8410), .S1(n7217), .Y(n7119) );
  OA22XL U10243 ( .A0(\xArray[14][44] ), .A1(n8270), .B0(\xArray[2][44] ), 
        .B1(n8185), .Y(n1375) );
  OA22XL U10244 ( .A0(\xArray[4][43] ), .A1(n8187), .B0(\xArray[0][43] ), .B1(
        n8258), .Y(n1078) );
  OA22XL U10245 ( .A0(\xArray[0][45] ), .A1(n8193), .B0(\xArray[12][45] ), 
        .B1(n8263), .Y(n1918) );
  OA22XL U10246 ( .A0(\xArray[15][45] ), .A1(n8193), .B0(\xArray[11][45] ), 
        .B1(n8263), .Y(n1917) );
  OA22XL U10247 ( .A0(\xArray[14][45] ), .A1(n8271), .B0(\xArray[2][45] ), 
        .B1(n8185), .Y(n1371) );
  OA22XL U10248 ( .A0(\xArray[0][46] ), .A1(n8193), .B0(\xArray[12][46] ), 
        .B1(n8263), .Y(n1909) );
  OA22XL U10249 ( .A0(\xArray[4][44] ), .A1(n6707), .B0(\xArray[0][44] ), .B1(
        n8254), .Y(n1073) );
  OA22XL U10250 ( .A0(\xArray[5][42] ), .A1(n8194), .B0(\xArray[1][42] ), .B1(
        n8255), .Y(n849) );
  OA22XL U10251 ( .A0(\xArray[5][43] ), .A1(n8194), .B0(\xArray[1][43] ), .B1(
        n8264), .Y(n846) );
  OA22XL U10252 ( .A0(\xArray[5][44] ), .A1(n8194), .B0(\xArray[1][44] ), .B1(
        n8253), .Y(n843) );
  AOI2BB2XL U10253 ( .B0(n9022), .B1(n8207), .A0N(\xArray[10][47] ), .A1N(
        n8253), .Y(n1897) );
  AOI2BB2XL U10254 ( .B0(n9014), .B1(n8217), .A0N(\xArray[10][48] ), .A1N(
        n8253), .Y(n1888) );
  OA22XL U10255 ( .A0(\xArray[4][46] ), .A1(n6707), .B0(\xArray[0][46] ), .B1(
        n8258), .Y(n1063) );
  OA22XL U10256 ( .A0(\xArray[4][47] ), .A1(n8186), .B0(\xArray[0][47] ), .B1(
        n8254), .Y(n1058) );
  OA22XL U10257 ( .A0(\xArray[14][48] ), .A1(n8273), .B0(\xArray[2][48] ), 
        .B1(n8184), .Y(n1359) );
  OA22XL U10258 ( .A0(\xArray[14][49] ), .A1(n8272), .B0(\xArray[2][49] ), 
        .B1(n8184), .Y(n1355) );
  OA22XL U10259 ( .A0(\xArray[15][48] ), .A1(n8198), .B0(\xArray[11][48] ), 
        .B1(n8262), .Y(n1890) );
  OA22XL U10260 ( .A0(\xArray[15][49] ), .A1(n8193), .B0(\xArray[11][49] ), 
        .B1(n8262), .Y(n1881) );
  OA22XL U10261 ( .A0(\xArray[1][48] ), .A1(n8199), .B0(\xArray[13][48] ), 
        .B1(n8267), .Y(n1599) );
  OA22XL U10262 ( .A0(\xArray[1][49] ), .A1(n8199), .B0(\xArray[13][49] ), 
        .B1(n8267), .Y(n1596) );
  OA22XL U10263 ( .A0(n8313), .A1(n1386), .B0(n7730), .B1(n1619), .Y(n1946) );
  OA22XL U10264 ( .A0(n8313), .A1(n1390), .B0(n7730), .B1(n1622), .Y(n1955) );
  MX4XL U10265 ( .A(\bArray[12][44] ), .B(\bArray[13][44] ), .C(
        \bArray[14][44] ), .D(\bArray[15][44] ), .S0(n8410), .S1(n7212), .Y(
        n7120) );
  MX4XL U10266 ( .A(\bArray[8][44] ), .B(\bArray[9][44] ), .C(\bArray[10][44] ), .D(\bArray[11][44] ), .S0(n7210), .S1(n7222), .Y(n7121) );
  AOI2BB2XL U10267 ( .B0(n9024), .B1(n8217), .A0N(\xArray[15][46] ), .A1N(
        n8257), .Y(n1064) );
  AOI2BB2XL U10268 ( .B0(n9016), .B1(n8217), .A0N(\xArray[15][47] ), .A1N(
        n8257), .Y(n1059) );
  INVXL U10269 ( .A(\xArray[5][35] ), .Y(n9114) );
  INVXL U10270 ( .A(\xArray[5][36] ), .Y(n9106) );
  NAND2BX1 U10271 ( .AN(n440), .B(n441), .Y(N34067) );
  NAND2BX1 U10272 ( .AN(n448), .B(n449), .Y(N34066) );
  INVXL U10273 ( .A(\xArray[9][35] ), .Y(n9116) );
  INVXL U10274 ( .A(\xArray[9][36] ), .Y(n9108) );
  INVXL U10275 ( .A(\xArray[6][35] ), .Y(n9115) );
  INVXL U10276 ( .A(\xArray[6][34] ), .Y(n9123) );
  INVXL U10277 ( .A(\xArray[10][35] ), .Y(n9117) );
  INVXL U10278 ( .A(\xArray[10][34] ), .Y(n9125) );
  OA22XL U10279 ( .A0(\xArray[0][48] ), .A1(n8194), .B0(\xArray[12][48] ), 
        .B1(n8263), .Y(n1891) );
  OA22XL U10280 ( .A0(\xArray[0][49] ), .A1(n8200), .B0(\xArray[12][49] ), 
        .B1(n8262), .Y(n1882) );
  OA22XL U10281 ( .A0(\xArray[5][45] ), .A1(n8194), .B0(\xArray[1][45] ), .B1(
        n8253), .Y(n840) );
  OA22XL U10282 ( .A0(\xArray[5][46] ), .A1(n8194), .B0(\xArray[1][46] ), .B1(
        n8253), .Y(n837) );
  AOI2BB2XL U10283 ( .B0(n9006), .B1(n8216), .A0N(\xArray[10][49] ), .A1N(
        n8253), .Y(n1879) );
  AOI2BB2XL U10284 ( .B0(n8998), .B1(n8207), .A0N(\xArray[10][50] ), .A1N(
        n8253), .Y(n1870) );
  OA22XL U10285 ( .A0(\xArray[4][48] ), .A1(n8198), .B0(\xArray[0][48] ), .B1(
        n8258), .Y(n1053) );
  OA22XL U10286 ( .A0(\xArray[4][49] ), .A1(n8198), .B0(\xArray[0][49] ), .B1(
        n8254), .Y(n1048) );
  OA22XL U10287 ( .A0(\xArray[14][50] ), .A1(n8273), .B0(\xArray[2][50] ), 
        .B1(n8184), .Y(n1351) );
  OA22XL U10288 ( .A0(\xArray[14][51] ), .A1(n8272), .B0(\xArray[2][51] ), 
        .B1(n8184), .Y(n1347) );
  OA22XL U10289 ( .A0(\xArray[15][50] ), .A1(n8200), .B0(\xArray[11][50] ), 
        .B1(n8262), .Y(n1872) );
  OA22XL U10290 ( .A0(\xArray[15][51] ), .A1(n8200), .B0(\xArray[11][51] ), 
        .B1(n8262), .Y(n1863) );
  OA22XL U10291 ( .A0(\xArray[1][50] ), .A1(n8199), .B0(\xArray[13][50] ), 
        .B1(n8267), .Y(n1593) );
  OA22XL U10292 ( .A0(\xArray[1][51] ), .A1(n8199), .B0(\xArray[13][51] ), 
        .B1(n8267), .Y(n1590) );
  OA22XL U10293 ( .A0(n8313), .A1(n1382), .B0(n7730), .B1(n1616), .Y(n1937) );
  OA22XL U10294 ( .A0(n8323), .A1(n1378), .B0(n7730), .B1(n1613), .Y(n1928) );
  AOI2BB2XL U10295 ( .B0(n9008), .B1(n8217), .A0N(\xArray[15][48] ), .A1N(
        n8257), .Y(n1054) );
  AOI2BB2XL U10296 ( .B0(n9000), .B1(n8217), .A0N(\xArray[15][49] ), .A1N(
        n8257), .Y(n1049) );
  INVXL U10297 ( .A(\xArray[5][37] ), .Y(n9098) );
  NAND2BX1 U10298 ( .AN(n424), .B(n425), .Y(N34069) );
  NAND2BX1 U10299 ( .AN(n432), .B(n433), .Y(N34068) );
  INVXL U10300 ( .A(\xArray[9][37] ), .Y(n9100) );
  INVXL U10301 ( .A(\xArray[6][37] ), .Y(n9099) );
  INVXL U10302 ( .A(\xArray[6][36] ), .Y(n9107) );
  INVXL U10303 ( .A(\xArray[10][37] ), .Y(n9101) );
  INVXL U10304 ( .A(\xArray[10][36] ), .Y(n9109) );
  OA22XL U10305 ( .A0(\xArray[0][50] ), .A1(n8200), .B0(\xArray[12][50] ), 
        .B1(n8262), .Y(n1873) );
  OA22XL U10306 ( .A0(\xArray[0][51] ), .A1(n8200), .B0(\xArray[12][51] ), 
        .B1(n8262), .Y(n1864) );
  OA22XL U10307 ( .A0(\xArray[5][47] ), .A1(n8194), .B0(\xArray[1][47] ), .B1(
        n8259), .Y(n834) );
  OA22XL U10308 ( .A0(\xArray[5][48] ), .A1(n8194), .B0(\xArray[1][48] ), .B1(
        n8259), .Y(n831) );
  AOI2BB2XL U10309 ( .B0(n8990), .B1(n8208), .A0N(\xArray[10][51] ), .A1N(
        n8253), .Y(n1861) );
  OA22XL U10310 ( .A0(\xArray[0][53] ), .A1(n8191), .B0(\xArray[12][53] ), 
        .B1(n8262), .Y(n1846) );
  AOI2BB2XL U10311 ( .B0(n8984), .B1(n8214), .A0N(\xArray[15][51] ), .A1N(
        n8259), .Y(n1039) );
  OA22XL U10312 ( .A0(\xArray[4][50] ), .A1(n6707), .B0(\xArray[0][50] ), .B1(
        n8258), .Y(n1043) );
  OA22XL U10313 ( .A0(\xArray[4][51] ), .A1(n8198), .B0(\xArray[0][51] ), .B1(
        n8254), .Y(n1038) );
  OA22XL U10314 ( .A0(\xArray[14][52] ), .A1(n8273), .B0(\xArray[2][52] ), 
        .B1(n8184), .Y(n1343) );
  OA22XL U10315 ( .A0(\xArray[14][53] ), .A1(n8272), .B0(\xArray[2][53] ), 
        .B1(n8184), .Y(n1339) );
  OA22XL U10316 ( .A0(\xArray[15][52] ), .A1(n8185), .B0(\xArray[11][52] ), 
        .B1(n8262), .Y(n1854) );
  OA22XL U10317 ( .A0(\xArray[15][53] ), .A1(n8195), .B0(\xArray[11][53] ), 
        .B1(n8262), .Y(n1845) );
  OA22XL U10318 ( .A0(\xArray[1][53] ), .A1(n8199), .B0(\xArray[13][53] ), 
        .B1(n8267), .Y(n1584) );
  OA22XL U10319 ( .A0(n8316), .A1(n1374), .B0(n7730), .B1(n1610), .Y(n1919) );
  OA22XL U10320 ( .A0(n8316), .A1(n1370), .B0(n7711), .B1(n1607), .Y(n1910) );
  AOI2BB2XL U10321 ( .B0(n8992), .B1(n8217), .A0N(\xArray[15][50] ), .A1N(
        n8257), .Y(n1044) );
  INVXL U10322 ( .A(\xArray[5][38] ), .Y(n9090) );
  INVXL U10323 ( .A(\xArray[5][39] ), .Y(n9082) );
  NAND2BX1 U10324 ( .AN(n408), .B(n409), .Y(N34071) );
  NAND2BX1 U10325 ( .AN(n416), .B(n417), .Y(N34070) );
  INVXL U10326 ( .A(\xArray[9][38] ), .Y(n9092) );
  INVXL U10327 ( .A(\xArray[9][39] ), .Y(n9084) );
  INVXL U10328 ( .A(\xArray[6][38] ), .Y(n9091) );
  INVXL U10329 ( .A(\xArray[10][39] ), .Y(n9085) );
  INVXL U10330 ( .A(\xArray[10][38] ), .Y(n9093) );
  OA22XL U10331 ( .A0(\xArray[1][52] ), .A1(n8199), .B0(\xArray[13][52] ), 
        .B1(n8267), .Y(n1587) );
  OA22XL U10332 ( .A0(\xArray[0][52] ), .A1(n8197), .B0(\xArray[12][52] ), 
        .B1(n8262), .Y(n1855) );
  OA22XL U10333 ( .A0(\xArray[5][49] ), .A1(n8194), .B0(\xArray[1][49] ), .B1(
        n8263), .Y(n828) );
  OA22XL U10334 ( .A0(\xArray[5][50] ), .A1(n8194), .B0(\xArray[1][50] ), .B1(
        n8263), .Y(n825) );
  AOI2BB2XL U10335 ( .B0(n8982), .B1(n8216), .A0N(\xArray[10][52] ), .A1N(
        n8253), .Y(n1852) );
  OA22XL U10336 ( .A0(\xArray[5][52] ), .A1(n8194), .B0(\xArray[1][52] ), .B1(
        n8254), .Y(n819) );
  AOI2BB2XL U10337 ( .B0(n8974), .B1(n8203), .A0N(\xArray[10][53] ), .A1N(
        n8253), .Y(n1843) );
  AOI2BB2XL U10338 ( .B0(n8966), .B1(n8203), .A0N(\xArray[10][54] ), .A1N(
        n8253), .Y(n1834) );
  OA22XL U10339 ( .A0(\xArray[0][54] ), .A1(n8184), .B0(\xArray[12][54] ), 
        .B1(n8262), .Y(n1837) );
  OA22XL U10340 ( .A0(\xArray[0][55] ), .A1(n8190), .B0(\xArray[12][55] ), 
        .B1(n8262), .Y(n1828) );
  AOI2BB2XL U10341 ( .B0(n8976), .B1(n8208), .A0N(\xArray[15][52] ), .A1N(
        n8259), .Y(n1034) );
  AOI2BB2XL U10342 ( .B0(n8968), .B1(n8214), .A0N(\xArray[15][53] ), .A1N(
        n8259), .Y(n1029) );
  OA22XL U10343 ( .A0(\xArray[4][52] ), .A1(n8192), .B0(\xArray[0][52] ), .B1(
        n8258), .Y(n1033) );
  OA22XL U10344 ( .A0(\xArray[4][53] ), .A1(n6707), .B0(\xArray[0][53] ), .B1(
        n8254), .Y(n1028) );
  OA22XL U10345 ( .A0(\xArray[14][54] ), .A1(n8273), .B0(\xArray[2][54] ), 
        .B1(n8184), .Y(n1335) );
  OA22XL U10346 ( .A0(\xArray[15][54] ), .A1(n8188), .B0(\xArray[11][54] ), 
        .B1(n8262), .Y(n1836) );
  OA22XL U10347 ( .A0(\xArray[1][54] ), .A1(n8199), .B0(\xArray[13][54] ), 
        .B1(n8267), .Y(n1581) );
  OA22XL U10348 ( .A0(\xArray[1][55] ), .A1(n8199), .B0(\xArray[13][55] ), 
        .B1(n8267), .Y(n1578) );
  OA22XL U10349 ( .A0(n8316), .A1(n1366), .B0(n7713), .B1(n1604), .Y(n1901) );
  MX4XL U10350 ( .A(\bArray[8][19] ), .B(\bArray[9][19] ), .C(\bArray[10][19] ), .D(\bArray[11][19] ), .S0(n6983), .S1(n6998), .Y(n6798) );
  MX4XL U10351 ( .A(\bArray[0][19] ), .B(\bArray[1][19] ), .C(\bArray[2][19] ), 
        .D(\bArray[3][19] ), .S0(n6983), .S1(n6998), .Y(n6800) );
  MX4XL U10352 ( .A(\bArray[12][19] ), .B(\bArray[13][19] ), .C(
        \bArray[14][19] ), .D(\bArray[15][19] ), .S0(n6983), .S1(n6998), .Y(
        n6797) );
  MX4XL U10353 ( .A(\bArray[8][18] ), .B(\bArray[9][18] ), .C(\bArray[10][18] ), .D(\bArray[11][18] ), .S0(n6982), .S1(n6997), .Y(n6794) );
  MX4XL U10354 ( .A(\bArray[12][18] ), .B(\bArray[13][18] ), .C(
        \bArray[14][18] ), .D(\bArray[15][18] ), .S0(n6982), .S1(n6997), .Y(
        n6793) );
  MX4XL U10355 ( .A(\bArray[0][18] ), .B(\bArray[1][18] ), .C(\bArray[2][18] ), 
        .D(\bArray[3][18] ), .S0(n6983), .S1(n6998), .Y(n6796) );
  INVXL U10356 ( .A(\xArray[5][40] ), .Y(n9074) );
  INVXL U10357 ( .A(\xArray[5][41] ), .Y(n9066) );
  NAND2BX1 U10358 ( .AN(n392), .B(n393), .Y(N34073) );
  NAND2BX1 U10359 ( .AN(n400), .B(n401), .Y(N34072) );
  INVXL U10360 ( .A(\xArray[9][40] ), .Y(n9076) );
  INVXL U10361 ( .A(\xArray[9][41] ), .Y(n9068) );
  INVXL U10362 ( .A(\xArray[6][40] ), .Y(n9075) );
  INVXL U10363 ( .A(\xArray[6][39] ), .Y(n9083) );
  INVXL U10364 ( .A(\xArray[10][40] ), .Y(n9077) );
  OA22XL U10365 ( .A0(\xArray[15][55] ), .A1(n8184), .B0(\xArray[11][55] ), 
        .B1(n8261), .Y(n1827) );
  OA22XL U10366 ( .A0(\xArray[14][55] ), .A1(n8273), .B0(\xArray[2][55] ), 
        .B1(n8184), .Y(n1331) );
  MX4XL U10367 ( .A(\bArray[4][19] ), .B(\bArray[5][19] ), .C(\bArray[6][19] ), 
        .D(\bArray[7][19] ), .S0(n6983), .S1(n6998), .Y(n6799) );
  MX4XL U10368 ( .A(\bArray[4][18] ), .B(\bArray[5][18] ), .C(\bArray[6][18] ), 
        .D(\bArray[7][18] ), .S0(n6983), .S1(n6998), .Y(n6795) );
  MX4XL U10369 ( .A(\bArray[8][17] ), .B(\bArray[9][17] ), .C(\bArray[10][17] ), .D(\bArray[11][17] ), .S0(n6982), .S1(n6997), .Y(n6790) );
  MX4XL U10370 ( .A(\bArray[0][17] ), .B(\bArray[1][17] ), .C(\bArray[2][17] ), 
        .D(\bArray[3][17] ), .S0(n6982), .S1(n6997), .Y(n6792) );
  MX4XL U10371 ( .A(\bArray[12][17] ), .B(\bArray[13][17] ), .C(
        \bArray[14][17] ), .D(\bArray[15][17] ), .S0(n6982), .S1(n6997), .Y(
        n6789) );
  MX4XL U10372 ( .A(\bArray[8][16] ), .B(\bArray[9][16] ), .C(\bArray[10][16] ), .D(\bArray[11][16] ), .S0(n6982), .S1(n6997), .Y(n6786) );
  MX4XL U10373 ( .A(\bArray[0][16] ), .B(\bArray[1][16] ), .C(\bArray[2][16] ), 
        .D(\bArray[3][16] ), .S0(n6982), .S1(n6997), .Y(n6788) );
  MX4XL U10374 ( .A(\bArray[12][16] ), .B(\bArray[13][16] ), .C(
        \bArray[14][16] ), .D(\bArray[15][16] ), .S0(n6982), .S1(n6997), .Y(
        n6785) );
  MX4XL U10375 ( .A(\bArray[4][17] ), .B(\bArray[5][17] ), .C(\bArray[6][17] ), 
        .D(\bArray[7][17] ), .S0(n6982), .S1(n6997), .Y(n6791) );
  MX4XL U10376 ( .A(\bArray[4][16] ), .B(\bArray[5][16] ), .C(\bArray[6][16] ), 
        .D(\bArray[7][16] ), .S0(n6982), .S1(n6997), .Y(n6787) );
  OA22XL U10377 ( .A0(\xArray[5][51] ), .A1(n8194), .B0(\xArray[1][51] ), .B1(
        n8263), .Y(n822) );
  OA22XL U10378 ( .A0(\xArray[5][53] ), .A1(n8194), .B0(\xArray[1][53] ), .B1(
        n8254), .Y(n816) );
  OA22XL U10379 ( .A0(\xArray[5][54] ), .A1(n8194), .B0(\xArray[1][54] ), .B1(
        n8254), .Y(n813) );
  AOI2BB2XL U10380 ( .B0(n8958), .B1(n8203), .A0N(\xArray[10][55] ), .A1N(
        n8253), .Y(n1825) );
  AOI2BB2XL U10381 ( .B0(n8950), .B1(n8209), .A0N(\xArray[10][56] ), .A1N(
        n8253), .Y(n1816) );
  OA22XL U10382 ( .A0(\xArray[0][56] ), .A1(n8187), .B0(\xArray[12][56] ), 
        .B1(n8261), .Y(n1819) );
  OA22XL U10383 ( .A0(\xArray[0][57] ), .A1(n8189), .B0(\xArray[12][57] ), 
        .B1(n8261), .Y(n1810) );
  AOI2BB2XL U10384 ( .B0(n8960), .B1(n8203), .A0N(\xArray[15][54] ), .A1N(
        n8259), .Y(n1024) );
  AOI2BB2XL U10385 ( .B0(n8952), .B1(n8203), .A0N(\xArray[15][55] ), .A1N(
        n8259), .Y(n1019) );
  OA22XL U10386 ( .A0(\xArray[4][54] ), .A1(n6707), .B0(\xArray[0][54] ), .B1(
        n8268), .Y(n1023) );
  OA22XL U10387 ( .A0(\xArray[4][55] ), .A1(n786), .B0(\xArray[0][55] ), .B1(
        n8268), .Y(n1018) );
  OA22XL U10388 ( .A0(\xArray[1][56] ), .A1(n8199), .B0(\xArray[13][56] ), 
        .B1(n8267), .Y(n1575) );
  OA22XL U10389 ( .A0(\xArray[1][57] ), .A1(n8199), .B0(\xArray[13][57] ), 
        .B1(n8267), .Y(n1572) );
  NAND2BX1 U10390 ( .AN(n376), .B(n377), .Y(N34075) );
  NAND2BX1 U10391 ( .AN(n384), .B(n385), .Y(N34074) );
  INVXL U10392 ( .A(\xArray[6][41] ), .Y(n9067) );
  INVXL U10393 ( .A(\xArray[10][41] ), .Y(n9069) );
  OA22XL U10394 ( .A0(\xArray[15][56] ), .A1(n8189), .B0(\xArray[11][56] ), 
        .B1(n8261), .Y(n1818) );
  OA22XL U10395 ( .A0(\xArray[15][57] ), .A1(n8189), .B0(\xArray[11][57] ), 
        .B1(n8261), .Y(n1809) );
  OA22XL U10396 ( .A0(\xArray[14][56] ), .A1(n8273), .B0(\xArray[2][56] ), 
        .B1(n8184), .Y(n1327) );
  AOI2BB2XL U10397 ( .B0(n8942), .B1(n8214), .A0N(\xArray[10][57] ), .A1N(
        n8253), .Y(n1807) );
  OA22XL U10398 ( .A0(\xArray[0][58] ), .A1(n8189), .B0(\xArray[12][58] ), 
        .B1(n8261), .Y(n1801) );
  OA22XL U10399 ( .A0(\xArray[0][59] ), .A1(n8189), .B0(\xArray[12][59] ), 
        .B1(n8261), .Y(n1792) );
  OA22XL U10400 ( .A0(\xArray[4][56] ), .A1(n786), .B0(\xArray[0][56] ), .B1(
        n8268), .Y(n1013) );
  OA22XL U10401 ( .A0(\xArray[4][57] ), .A1(n786), .B0(\xArray[0][57] ), .B1(
        n8268), .Y(n1008) );
  OA22XL U10402 ( .A0(\xArray[1][58] ), .A1(n8199), .B0(\xArray[13][58] ), 
        .B1(n8267), .Y(n1569) );
  OA22XL U10403 ( .A0(n8321), .A1(n1346), .B0(n7711), .B1(n1589), .Y(n1856) );
  MX4XL U10404 ( .A(\bArray[8][23] ), .B(\bArray[9][23] ), .C(\bArray[10][23] ), .D(\bArray[11][23] ), .S0(n6984), .S1(n6999), .Y(n6814) );
  MX4XL U10405 ( .A(\bArray[0][23] ), .B(\bArray[1][23] ), .C(\bArray[2][23] ), 
        .D(\bArray[3][23] ), .S0(n6984), .S1(n6999), .Y(n6816) );
  MX4XL U10406 ( .A(\bArray[12][23] ), .B(\bArray[13][23] ), .C(
        \bArray[14][23] ), .D(\bArray[15][23] ), .S0(n6984), .S1(n6999), .Y(
        n6813) );
  MX4XL U10407 ( .A(\bArray[8][22] ), .B(\bArray[9][22] ), .C(\bArray[10][22] ), .D(\bArray[11][22] ), .S0(n6984), .S1(n6999), .Y(n6810) );
  MX4XL U10408 ( .A(\bArray[0][22] ), .B(\bArray[1][22] ), .C(\bArray[2][22] ), 
        .D(\bArray[3][22] ), .S0(n6984), .S1(n6999), .Y(n6812) );
  MX4XL U10409 ( .A(\bArray[12][22] ), .B(\bArray[13][22] ), .C(
        \bArray[14][22] ), .D(\bArray[15][22] ), .S0(n6984), .S1(n6999), .Y(
        n6809) );
  MX4XL U10410 ( .A(\bArray[8][21] ), .B(\bArray[9][21] ), .C(\bArray[10][21] ), .D(\bArray[11][21] ), .S0(n6983), .S1(n6998), .Y(n6806) );
  MX4XL U10411 ( .A(\bArray[0][21] ), .B(\bArray[1][21] ), .C(\bArray[2][21] ), 
        .D(\bArray[3][21] ), .S0(n6984), .S1(n6999), .Y(n6808) );
  MX4XL U10412 ( .A(\bArray[12][21] ), .B(\bArray[13][21] ), .C(
        \bArray[14][21] ), .D(\bArray[15][21] ), .S0(n6983), .S1(n6998), .Y(
        n6805) );
  MX4XL U10413 ( .A(\bArray[8][20] ), .B(\bArray[9][20] ), .C(\bArray[10][20] ), .D(\bArray[11][20] ), .S0(n6983), .S1(n6998), .Y(n6802) );
  MX4XL U10414 ( .A(\bArray[0][20] ), .B(\bArray[1][20] ), .C(\bArray[2][20] ), 
        .D(\bArray[3][20] ), .S0(n6983), .S1(n6998), .Y(n6804) );
  MX4XL U10415 ( .A(\bArray[12][20] ), .B(\bArray[13][20] ), .C(
        \bArray[14][20] ), .D(\bArray[15][20] ), .S0(n6983), .S1(n6998), .Y(
        n6801) );
  NAND2BX1 U10416 ( .AN(n368), .B(n369), .Y(N34076) );
  OA22XL U10417 ( .A0(\xArray[15][58] ), .A1(n8189), .B0(\xArray[11][58] ), 
        .B1(n8261), .Y(n1800) );
  OA22XL U10418 ( .A0(\xArray[15][59] ), .A1(n8189), .B0(\xArray[11][59] ), 
        .B1(n8261), .Y(n1791) );
  OA22XL U10419 ( .A0(\xArray[14][57] ), .A1(n8273), .B0(\xArray[2][57] ), 
        .B1(n8184), .Y(n1323) );
  OA22XL U10420 ( .A0(\xArray[14][58] ), .A1(n8273), .B0(\xArray[2][58] ), 
        .B1(n8184), .Y(n1319) );
  MX4XL U10421 ( .A(\bArray[4][23] ), .B(\bArray[5][23] ), .C(\bArray[6][23] ), 
        .D(\bArray[7][23] ), .S0(n6984), .S1(n6999), .Y(n6815) );
  MX4XL U10422 ( .A(\bArray[4][22] ), .B(\bArray[5][22] ), .C(\bArray[6][22] ), 
        .D(\bArray[7][22] ), .S0(n6984), .S1(n6999), .Y(n6811) );
  MX4XL U10423 ( .A(\bArray[4][21] ), .B(\bArray[5][21] ), .C(\bArray[6][21] ), 
        .D(\bArray[7][21] ), .S0(n6983), .S1(n6998), .Y(n6807) );
  MX4XL U10424 ( .A(\bArray[4][20] ), .B(\bArray[5][20] ), .C(\bArray[6][20] ), 
        .D(\bArray[7][20] ), .S0(n6983), .S1(n6998), .Y(n6803) );
  AOI2BB2XL U10425 ( .B0(n8934), .B1(n8214), .A0N(\xArray[10][58] ), .A1N(
        n8253), .Y(n1798) );
  AOI2BB2XL U10426 ( .B0(n8926), .B1(n8208), .A0N(\xArray[10][59] ), .A1N(
        n8253), .Y(n1789) );
  OA22XL U10427 ( .A0(\xArray[0][60] ), .A1(n8189), .B0(\xArray[12][60] ), 
        .B1(n8261), .Y(n1783) );
  AOI2BB2XL U10428 ( .B0(n8920), .B1(n8214), .A0N(\xArray[15][59] ), .A1N(
        n8258), .Y(n999) );
  OA22XL U10429 ( .A0(\xArray[4][58] ), .A1(n786), .B0(\xArray[0][58] ), .B1(
        n8268), .Y(n1003) );
  OA22XL U10430 ( .A0(\xArray[4][59] ), .A1(n8196), .B0(\xArray[0][59] ), .B1(
        n8268), .Y(n998) );
  OA22XL U10431 ( .A0(n8321), .A1(n1338), .B0(n7726), .B1(n1583), .Y(n1838) );
  OA22XL U10432 ( .A0(n8321), .A1(n1342), .B0(n7711), .B1(n1586), .Y(n1847) );
  NAND2BX1 U10433 ( .AN(n352), .B(n353), .Y(N34078) );
  NAND2BX1 U10434 ( .AN(n360), .B(n361), .Y(N34077) );
  OA22XL U10435 ( .A0(\xArray[15][60] ), .A1(n8188), .B0(\xArray[11][60] ), 
        .B1(n8261), .Y(n1782) );
  OA22XL U10436 ( .A0(\xArray[14][59] ), .A1(n8273), .B0(\xArray[2][59] ), 
        .B1(n8184), .Y(n1315) );
  OA22XL U10437 ( .A0(\xArray[14][60] ), .A1(n8273), .B0(\xArray[2][60] ), 
        .B1(n8184), .Y(n1311) );
  OA22XL U10438 ( .A0(\xArray[0][61] ), .A1(n8188), .B0(\xArray[12][61] ), 
        .B1(n8260), .Y(n1774) );
  AOI2BB2XL U10439 ( .B0(n8912), .B1(n8213), .A0N(\xArray[15][60] ), .A1N(
        n8257), .Y(n994) );
  OA22XL U10440 ( .A0(\xArray[14][61] ), .A1(n8273), .B0(\xArray[2][61] ), 
        .B1(n8184), .Y(n1307) );
  OA22XL U10441 ( .A0(n8321), .A1(n1334), .B0(n7711), .B1(n1580), .Y(n1829) );
  OA22XL U10442 ( .A0(n8321), .A1(n1330), .B0(n7726), .B1(n1577), .Y(n1820) );
  OA22XL U10443 ( .A0(\xArray[4][60] ), .A1(n8196), .B0(\xArray[0][60] ), .B1(
        n8268), .Y(n993) );
  MX4XL U10444 ( .A(\bArray[8][27] ), .B(\bArray[9][27] ), .C(\bArray[10][27] ), .D(\bArray[11][27] ), .S0(n6985), .S1(n8413), .Y(n6830) );
  MX4XL U10445 ( .A(\bArray[0][27] ), .B(\bArray[1][27] ), .C(\bArray[2][27] ), 
        .D(\bArray[3][27] ), .S0(n6985), .S1(n8413), .Y(n6832) );
  MX4XL U10446 ( .A(\bArray[12][27] ), .B(\bArray[13][27] ), .C(
        \bArray[14][27] ), .D(\bArray[15][27] ), .S0(n6985), .S1(n8413), .Y(
        n6829) );
  MX4XL U10447 ( .A(\bArray[8][26] ), .B(\bArray[9][26] ), .C(\bArray[10][26] ), .D(\bArray[11][26] ), .S0(n6985), .S1(n8413), .Y(n6826) );
  MX4XL U10448 ( .A(\bArray[0][26] ), .B(\bArray[1][26] ), .C(\bArray[2][26] ), 
        .D(\bArray[3][26] ), .S0(n6985), .S1(n8413), .Y(n6828) );
  MX4XL U10449 ( .A(\bArray[12][26] ), .B(\bArray[13][26] ), .C(
        \bArray[14][26] ), .D(\bArray[15][26] ), .S0(n6985), .S1(n8413), .Y(
        n6825) );
  MX4XL U10450 ( .A(\bArray[8][25] ), .B(\bArray[9][25] ), .C(\bArray[10][25] ), .D(\bArray[11][25] ), .S0(n6985), .S1(n6997), .Y(n6822) );
  MX4XL U10451 ( .A(\bArray[0][25] ), .B(\bArray[1][25] ), .C(\bArray[2][25] ), 
        .D(\bArray[3][25] ), .S0(n6985), .S1(n8413), .Y(n6824) );
  MX4XL U10452 ( .A(\bArray[12][25] ), .B(\bArray[13][25] ), .C(
        \bArray[14][25] ), .D(\bArray[15][25] ), .S0(n6985), .S1(n6999), .Y(
        n6821) );
  MX4XL U10453 ( .A(\bArray[8][24] ), .B(\bArray[9][24] ), .C(\bArray[10][24] ), .D(\bArray[11][24] ), .S0(n6984), .S1(n6999), .Y(n6818) );
  MX4XL U10454 ( .A(\bArray[0][24] ), .B(\bArray[1][24] ), .C(\bArray[2][24] ), 
        .D(\bArray[3][24] ), .S0(n6984), .S1(n6999), .Y(n6820) );
  MX4XL U10455 ( .A(\bArray[12][24] ), .B(\bArray[13][24] ), .C(
        \bArray[14][24] ), .D(\bArray[15][24] ), .S0(n6984), .S1(n6999), .Y(
        n6817) );
  NAND2BX1 U10456 ( .AN(n336), .B(n337), .Y(N34080) );
  NAND2BX1 U10457 ( .AN(n344), .B(n345), .Y(N34079) );
  OA22XL U10458 ( .A0(\xArray[15][61] ), .A1(n8188), .B0(\xArray[11][61] ), 
        .B1(n8260), .Y(n1773) );
  MX4XL U10459 ( .A(\bArray[4][27] ), .B(\bArray[5][27] ), .C(\bArray[6][27] ), 
        .D(\bArray[7][27] ), .S0(n6985), .S1(n8413), .Y(n6831) );
  MX4XL U10460 ( .A(\bArray[4][26] ), .B(\bArray[5][26] ), .C(\bArray[6][26] ), 
        .D(\bArray[7][26] ), .S0(n6985), .S1(n8413), .Y(n6827) );
  MX4XL U10461 ( .A(\bArray[4][25] ), .B(\bArray[5][25] ), .C(\bArray[6][25] ), 
        .D(\bArray[7][25] ), .S0(n6985), .S1(n6995), .Y(n6823) );
  MX4XL U10462 ( .A(\bArray[4][24] ), .B(\bArray[5][24] ), .C(\bArray[6][24] ), 
        .D(\bArray[7][24] ), .S0(n6984), .S1(n6999), .Y(n6819) );
  OA22XL U10463 ( .A0(\xArray[0][62] ), .A1(n8188), .B0(\xArray[12][62] ), 
        .B1(n8260), .Y(n1765) );
  AOI2BB2XL U10464 ( .B0(n8904), .B1(n8213), .A0N(\xArray[15][61] ), .A1N(
        n8258), .Y(n989) );
  OA22XL U10465 ( .A0(\xArray[4][61] ), .A1(n8196), .B0(\xArray[0][61] ), .B1(
        n8268), .Y(n988) );
  OA22XL U10466 ( .A0(\xArray[15][62] ), .A1(n8188), .B0(\xArray[11][62] ), 
        .B1(n8260), .Y(n1764) );
  OA22XL U10467 ( .A0(n8321), .A1(n1326), .B0(n7725), .B1(n1574), .Y(n1811) );
  NAND2BX1 U10468 ( .AN(n320), .B(n321), .Y(N34082) );
  NAND2BX1 U10469 ( .AN(n328), .B(n329), .Y(N34081) );
  OA22XL U10470 ( .A0(\xArray[14][62] ), .A1(n8273), .B0(\xArray[2][62] ), 
        .B1(n8184), .Y(n1303) );
  AOI2BB2XL U10471 ( .B0(n8902), .B1(n8210), .A0N(\xArray[10][62] ), .A1N(
        n8253), .Y(n1762) );
  AOI2BB2XL U10472 ( .B0(n8896), .B1(n8213), .A0N(\xArray[15][62] ), .A1N(
        n8258), .Y(n984) );
  OA22XL U10473 ( .A0(\xArray[4][62] ), .A1(n8196), .B0(\xArray[0][62] ), .B1(
        n8268), .Y(n983) );
  OA22XL U10474 ( .A0(n8321), .A1(n1322), .B0(n7729), .B1(n1571), .Y(n1802) );
  OA22XL U10475 ( .A0(n8321), .A1(n1318), .B0(n7726), .B1(n1568), .Y(n1793) );
  MX4XL U10476 ( .A(\bArray[8][31] ), .B(\bArray[9][31] ), .C(\bArray[10][31] ), .D(\bArray[11][31] ), .S0(n6986), .S1(N1758), .Y(n6846) );
  MX4XL U10477 ( .A(\bArray[0][31] ), .B(\bArray[1][31] ), .C(\bArray[2][31] ), 
        .D(\bArray[3][31] ), .S0(n6987), .S1(n7000), .Y(n6848) );
  MX4XL U10478 ( .A(\bArray[12][31] ), .B(\bArray[13][31] ), .C(
        \bArray[14][31] ), .D(\bArray[15][31] ), .S0(n6986), .S1(N1758), .Y(
        n6845) );
  MX4XL U10479 ( .A(\bArray[8][30] ), .B(\bArray[9][30] ), .C(\bArray[10][30] ), .D(\bArray[11][30] ), .S0(n6986), .S1(N1758), .Y(n6842) );
  MX4XL U10480 ( .A(\bArray[0][30] ), .B(\bArray[1][30] ), .C(\bArray[2][30] ), 
        .D(\bArray[3][30] ), .S0(n6986), .S1(N1758), .Y(n6844) );
  MX4XL U10481 ( .A(\bArray[12][30] ), .B(\bArray[13][30] ), .C(
        \bArray[14][30] ), .D(\bArray[15][30] ), .S0(n6986), .S1(n6997), .Y(
        n6841) );
  MX4XL U10482 ( .A(\bArray[8][29] ), .B(\bArray[9][29] ), .C(\bArray[10][29] ), .D(\bArray[11][29] ), .S0(n6986), .S1(n6999), .Y(n6838) );
  MX4XL U10483 ( .A(\bArray[0][29] ), .B(\bArray[1][29] ), .C(\bArray[2][29] ), 
        .D(\bArray[3][29] ), .S0(n6986), .S1(n6998), .Y(n6840) );
  MX4XL U10484 ( .A(\bArray[12][29] ), .B(\bArray[13][29] ), .C(
        \bArray[14][29] ), .D(\bArray[15][29] ), .S0(n6986), .S1(n6999), .Y(
        n6837) );
  MX4XL U10485 ( .A(\bArray[12][28] ), .B(\bArray[13][28] ), .C(
        \bArray[14][28] ), .D(\bArray[15][28] ), .S0(n6985), .S1(n8413), .Y(
        n6833) );
  MX4XL U10486 ( .A(\bArray[8][28] ), .B(\bArray[9][28] ), .C(\bArray[10][28] ), .D(\bArray[11][28] ), .S0(n6986), .S1(n6999), .Y(n6834) );
  MX4XL U10487 ( .A(\bArray[0][28] ), .B(\bArray[1][28] ), .C(\bArray[2][28] ), 
        .D(\bArray[3][28] ), .S0(n6986), .S1(n6995), .Y(n6836) );
  NAND2BX1 U10488 ( .AN(n304), .B(n305), .Y(N34084) );
  NAND2BX1 U10489 ( .AN(n312), .B(n313), .Y(N34083) );
  MX4XL U10490 ( .A(\bArray[4][31] ), .B(\bArray[5][31] ), .C(\bArray[6][31] ), 
        .D(\bArray[7][31] ), .S0(n6987), .S1(n7000), .Y(n6847) );
  MX4XL U10491 ( .A(\bArray[4][30] ), .B(\bArray[5][30] ), .C(\bArray[6][30] ), 
        .D(\bArray[7][30] ), .S0(n6986), .S1(n8413), .Y(n6843) );
  MX4XL U10492 ( .A(\bArray[4][29] ), .B(\bArray[5][29] ), .C(\bArray[6][29] ), 
        .D(\bArray[7][29] ), .S0(n6986), .S1(n6998), .Y(n6839) );
  MX4XL U10493 ( .A(\bArray[4][28] ), .B(\bArray[5][28] ), .C(\bArray[6][28] ), 
        .D(\bArray[7][28] ), .S0(n6986), .S1(n6994), .Y(n6835) );
  OA22XL U10494 ( .A0(\xArray[15][63] ), .A1(n8187), .B0(\xArray[11][63] ), 
        .B1(n8260), .Y(n1755) );
  OA22XL U10495 ( .A0(n8321), .A1(n1310), .B0(n7729), .B1(n1562), .Y(n1775) );
  OA22XL U10496 ( .A0(n8321), .A1(n1314), .B0(n7711), .B1(n1565), .Y(n1784) );
  NAND2BX1 U10497 ( .AN(n288), .B(n289), .Y(N34086) );
  NAND2BX1 U10498 ( .AN(n296), .B(n297), .Y(N34085) );
  OA22XL U10499 ( .A0(\xArray[0][63] ), .A1(n8187), .B0(\xArray[12][63] ), 
        .B1(n8260), .Y(n1756) );
  AOI2BB2XL U10500 ( .B0(n8888), .B1(n8213), .A0N(\xArray[15][63] ), .A1N(
        n8258), .Y(n979) );
  OA22XL U10501 ( .A0(\xArray[1][63] ), .A1(n8198), .B0(\xArray[13][63] ), 
        .B1(n8270), .Y(n1554) );
  OA22XL U10502 ( .A0(\xArray[4][63] ), .A1(n8196), .B0(\xArray[0][63] ), .B1(
        n8268), .Y(n978) );
  OA22XL U10503 ( .A0(n8321), .A1(n1306), .B0(n7720), .B1(n1559), .Y(n1766) );
  OA22XL U10504 ( .A0(n8321), .A1(n1302), .B0(n7720), .B1(n1556), .Y(n1757) );
  MX4XL U10505 ( .A(\bArray[8][35] ), .B(\bArray[9][35] ), .C(\bArray[10][35] ), .D(\bArray[11][35] ), .S0(n6988), .S1(n6998), .Y(n6862) );
  MX4XL U10506 ( .A(\bArray[0][35] ), .B(\bArray[1][35] ), .C(\bArray[2][35] ), 
        .D(\bArray[3][35] ), .S0(n6988), .S1(n7001), .Y(n6864) );
  MX4XL U10507 ( .A(\bArray[12][35] ), .B(\bArray[13][35] ), .C(
        \bArray[14][35] ), .D(\bArray[15][35] ), .S0(n6988), .S1(n6999), .Y(
        n6861) );
  MX4XL U10508 ( .A(\bArray[8][34] ), .B(\bArray[9][34] ), .C(\bArray[10][34] ), .D(\bArray[11][34] ), .S0(n6987), .S1(n7000), .Y(n6858) );
  MX4XL U10509 ( .A(\bArray[0][34] ), .B(\bArray[1][34] ), .C(\bArray[2][34] ), 
        .D(\bArray[3][34] ), .S0(n6988), .S1(n6993), .Y(n6860) );
  MX4XL U10510 ( .A(\bArray[12][34] ), .B(\bArray[13][34] ), .C(
        \bArray[14][34] ), .D(\bArray[15][34] ), .S0(n6987), .S1(n7000), .Y(
        n6857) );
  MX4XL U10511 ( .A(\bArray[8][33] ), .B(\bArray[9][33] ), .C(\bArray[10][33] ), .D(\bArray[11][33] ), .S0(n6987), .S1(n7000), .Y(n6854) );
  MX4XL U10512 ( .A(\bArray[0][33] ), .B(\bArray[1][33] ), .C(\bArray[2][33] ), 
        .D(\bArray[3][33] ), .S0(n6987), .S1(n7000), .Y(n6856) );
  MX4XL U10513 ( .A(\bArray[12][33] ), .B(\bArray[13][33] ), .C(
        \bArray[14][33] ), .D(\bArray[15][33] ), .S0(n6987), .S1(n7000), .Y(
        n6853) );
  MX4XL U10514 ( .A(\bArray[8][32] ), .B(\bArray[9][32] ), .C(\bArray[10][32] ), .D(\bArray[11][32] ), .S0(n6987), .S1(n7000), .Y(n6850) );
  MX4XL U10515 ( .A(\bArray[0][32] ), .B(\bArray[1][32] ), .C(\bArray[2][32] ), 
        .D(\bArray[3][32] ), .S0(n6987), .S1(n7000), .Y(n6852) );
  MX4XL U10516 ( .A(\bArray[12][32] ), .B(\bArray[13][32] ), .C(
        \bArray[14][32] ), .D(\bArray[15][32] ), .S0(n6987), .S1(n7000), .Y(
        n6849) );
  NAND2BX1 U10517 ( .AN(n280), .B(n281), .Y(N34087) );
  NAND2BX1 U10518 ( .AN(n272), .B(n273), .Y(N34088) );
  OA22XL U10519 ( .A0(\xArray[14][63] ), .A1(n8273), .B0(\xArray[2][63] ), 
        .B1(n8184), .Y(n1299) );
  MX4XL U10520 ( .A(\bArray[4][35] ), .B(\bArray[5][35] ), .C(\bArray[6][35] ), 
        .D(\bArray[7][35] ), .S0(n6988), .S1(n6997), .Y(n6863) );
  MX4XL U10521 ( .A(\bArray[4][34] ), .B(\bArray[5][34] ), .C(\bArray[6][34] ), 
        .D(\bArray[7][34] ), .S0(n6987), .S1(n7000), .Y(n6859) );
  MX4XL U10522 ( .A(\bArray[4][33] ), .B(\bArray[5][33] ), .C(\bArray[6][33] ), 
        .D(\bArray[7][33] ), .S0(n6987), .S1(n7000), .Y(n6855) );
  MX4XL U10523 ( .A(\bArray[4][32] ), .B(\bArray[5][32] ), .C(\bArray[6][32] ), 
        .D(\bArray[7][32] ), .S0(n6987), .S1(n7000), .Y(n6851) );
  OA22XL U10524 ( .A0(n8321), .A1(n1298), .B0(n7730), .B1(n1553), .Y(n1744) );
  NAND2BX1 U10525 ( .AN(n257), .B(n258), .Y(N34089) );
  OA22XL U10526 ( .A0(\xArray[5][63] ), .A1(n8189), .B0(\xArray[1][63] ), .B1(
        n8263), .Y(n785) );
  AOI2BB2XL U10527 ( .B0(n8894), .B1(n8210), .A0N(\xArray[10][63] ), .A1N(
        n8253), .Y(n1753) );
  MX4XL U10528 ( .A(\bArray[8][38] ), .B(\bArray[9][38] ), .C(\bArray[10][38] ), .D(\bArray[11][38] ), .S0(n6979), .S1(n6995), .Y(n6874) );
  MX4XL U10529 ( .A(\bArray[0][38] ), .B(\bArray[1][38] ), .C(\bArray[2][38] ), 
        .D(\bArray[3][38] ), .S0(n6979), .S1(N1758), .Y(n6876) );
  MX4XL U10530 ( .A(\bArray[12][38] ), .B(\bArray[13][38] ), .C(
        \bArray[14][38] ), .D(\bArray[15][38] ), .S0(n6982), .S1(n6993), .Y(
        n6873) );
  MX4XL U10531 ( .A(\bArray[8][37] ), .B(\bArray[9][37] ), .C(\bArray[10][37] ), .D(\bArray[11][37] ), .S0(n6988), .S1(n7001), .Y(n6870) );
  MX4XL U10532 ( .A(\bArray[0][37] ), .B(\bArray[1][37] ), .C(\bArray[2][37] ), 
        .D(\bArray[3][37] ), .S0(n6988), .S1(n7001), .Y(n6872) );
  MX4XL U10533 ( .A(\bArray[12][37] ), .B(\bArray[13][37] ), .C(
        \bArray[14][37] ), .D(\bArray[15][37] ), .S0(n6988), .S1(n7001), .Y(
        n6869) );
  MX4XL U10534 ( .A(\bArray[8][36] ), .B(\bArray[9][36] ), .C(\bArray[10][36] ), .D(\bArray[11][36] ), .S0(n6988), .S1(n7001), .Y(n6866) );
  MX4XL U10535 ( .A(\bArray[0][36] ), .B(\bArray[1][36] ), .C(\bArray[2][36] ), 
        .D(\bArray[3][36] ), .S0(n6988), .S1(n7001), .Y(n6868) );
  MX4XL U10536 ( .A(\bArray[12][36] ), .B(\bArray[13][36] ), .C(
        \bArray[14][36] ), .D(\bArray[15][36] ), .S0(n6988), .S1(n7001), .Y(
        n6865) );
  MX4XL U10537 ( .A(\bArray[4][38] ), .B(\bArray[5][38] ), .C(\bArray[6][38] ), 
        .D(\bArray[7][38] ), .S0(n6979), .S1(n6995), .Y(n6875) );
  MX4XL U10538 ( .A(\bArray[4][37] ), .B(\bArray[5][37] ), .C(\bArray[6][37] ), 
        .D(\bArray[7][37] ), .S0(n6988), .S1(n7001), .Y(n6871) );
  MX4XL U10539 ( .A(\bArray[4][36] ), .B(\bArray[5][36] ), .C(\bArray[6][36] ), 
        .D(\bArray[7][36] ), .S0(n6988), .S1(n7001), .Y(n6867) );
  NOR2BX1 U10540 ( .AN(n3638), .B(n5701), .Y(n3292) );
  NOR2BX1 U10541 ( .AN(n3078), .B(n5701), .Y(n2594) );
  NOR2X1 U10542 ( .A(n5703), .B(n5702), .Y(n3077) );
  CLKBUFX3 U10543 ( .A(N35189), .Y(n8404) );
  NAND2X1 U10544 ( .A(state[0]), .B(n6620), .Y(n241) );
  MX4XL U10545 ( .A(\xArray[0][2] ), .B(\xArray[1][2] ), .C(\xArray[2][2] ), 
        .D(\xArray[3][2] ), .S0(n7367), .S1(n8406), .Y(n7239) );
  MX4XL U10546 ( .A(\xArray[0][3] ), .B(\xArray[1][3] ), .C(\xArray[2][3] ), 
        .D(\xArray[3][3] ), .S0(n7367), .S1(n7361), .Y(n7243) );
  MX4XL U10547 ( .A(\xArray[0][4] ), .B(\xArray[1][4] ), .C(\xArray[2][4] ), 
        .D(\xArray[3][4] ), .S0(n7367), .S1(n7362), .Y(n7247) );
  MX4XL U10548 ( .A(\xArray[0][5] ), .B(\xArray[1][5] ), .C(\xArray[2][5] ), 
        .D(\xArray[3][5] ), .S0(n7367), .S1(n8406), .Y(n7251) );
  MX4XL U10549 ( .A(\xArray[0][6] ), .B(\xArray[1][6] ), .C(\xArray[2][6] ), 
        .D(\xArray[3][6] ), .S0(n7368), .S1(n7362), .Y(n7255) );
  MX4XL U10550 ( .A(\xArray[0][7] ), .B(\xArray[1][7] ), .C(\xArray[2][7] ), 
        .D(\xArray[3][7] ), .S0(n7368), .S1(n7363), .Y(n7259) );
  MX4XL U10551 ( .A(\xArray[0][8] ), .B(\xArray[1][8] ), .C(\xArray[2][8] ), 
        .D(\xArray[3][8] ), .S0(n7368), .S1(n7361), .Y(n7263) );
  MX4XL U10552 ( .A(\xArray[0][9] ), .B(\xArray[1][9] ), .C(\xArray[2][9] ), 
        .D(\xArray[3][9] ), .S0(n7369), .S1(n7361), .Y(n7267) );
  MX4XL U10553 ( .A(\xArray[0][10] ), .B(\xArray[1][10] ), .C(\xArray[2][10] ), 
        .D(\xArray[3][10] ), .S0(n7369), .S1(n7361), .Y(n7271) );
  MX4XL U10554 ( .A(\xArray[0][11] ), .B(\xArray[1][11] ), .C(\xArray[2][11] ), 
        .D(\xArray[3][11] ), .S0(n7369), .S1(n7361), .Y(n7275) );
  MX4XL U10555 ( .A(\xArray[0][12] ), .B(\xArray[1][12] ), .C(\xArray[2][12] ), 
        .D(\xArray[3][12] ), .S0(n7370), .S1(n7362), .Y(n7279) );
  MX4XL U10556 ( .A(\xArray[0][13] ), .B(\xArray[1][13] ), .C(\xArray[2][13] ), 
        .D(\xArray[3][13] ), .S0(n7370), .S1(n7362), .Y(n7283) );
  MX4XL U10557 ( .A(\xArray[0][14] ), .B(\xArray[1][14] ), .C(\xArray[2][14] ), 
        .D(\xArray[3][14] ), .S0(n7370), .S1(n7362), .Y(n7287) );
  MX4XL U10558 ( .A(\xArray[0][15] ), .B(\xArray[1][15] ), .C(\xArray[2][15] ), 
        .D(\xArray[3][15] ), .S0(n7371), .S1(n7363), .Y(n7291) );
  MX4XL U10559 ( .A(\xArray[0][16] ), .B(\xArray[1][16] ), .C(\xArray[2][16] ), 
        .D(\xArray[3][16] ), .S0(n7371), .S1(n7363), .Y(n7295) );
  MX4XL U10560 ( .A(\xArray[0][17] ), .B(\xArray[1][17] ), .C(\xArray[2][17] ), 
        .D(\xArray[3][17] ), .S0(n7371), .S1(n7363), .Y(n7299) );
  MX4XL U10561 ( .A(\xArray[0][18] ), .B(\xArray[1][18] ), .C(\xArray[2][18] ), 
        .D(\xArray[3][18] ), .S0(n7371), .S1(n7363), .Y(n7303) );
  MX4XL U10562 ( .A(\xArray[0][19] ), .B(\xArray[1][19] ), .C(\xArray[2][19] ), 
        .D(\xArray[3][19] ), .S0(n7372), .S1(n7364), .Y(n7307) );
  MX4XL U10563 ( .A(\xArray[0][20] ), .B(\xArray[1][20] ), .C(\xArray[2][20] ), 
        .D(\xArray[3][20] ), .S0(n7372), .S1(n7364), .Y(n7311) );
  MX4XL U10564 ( .A(\xArray[0][21] ), .B(\xArray[1][21] ), .C(\xArray[2][21] ), 
        .D(\xArray[3][21] ), .S0(n7372), .S1(n7364), .Y(n7315) );
  MX4XL U10565 ( .A(\xArray[0][22] ), .B(\xArray[1][22] ), .C(\xArray[2][22] ), 
        .D(\xArray[3][22] ), .S0(n7373), .S1(n7365), .Y(n7319) );
  MX4XL U10566 ( .A(\xArray[0][23] ), .B(\xArray[1][23] ), .C(\xArray[2][23] ), 
        .D(\xArray[3][23] ), .S0(n7373), .S1(n7365), .Y(n7323) );
  MX4XL U10567 ( .A(\xArray[0][24] ), .B(\xArray[1][24] ), .C(\xArray[2][24] ), 
        .D(\xArray[3][24] ), .S0(n7373), .S1(n7365), .Y(n7327) );
  MX4XL U10568 ( .A(\xArray[0][25] ), .B(\xArray[1][25] ), .C(\xArray[2][25] ), 
        .D(\xArray[3][25] ), .S0(n7373), .S1(n7366), .Y(n7331) );
  MX4XL U10569 ( .A(\xArray[0][26] ), .B(\xArray[1][26] ), .C(\xArray[2][26] ), 
        .D(\xArray[3][26] ), .S0(n7367), .S1(n7366), .Y(n7335) );
  MX4XL U10570 ( .A(\xArray[0][27] ), .B(\xArray[1][27] ), .C(\xArray[2][27] ), 
        .D(\xArray[3][27] ), .S0(n7370), .S1(n7366), .Y(n7339) );
  MX4XL U10571 ( .A(\xArray[0][28] ), .B(\xArray[1][28] ), .C(\xArray[2][28] ), 
        .D(\xArray[3][28] ), .S0(n7368), .S1(n7366), .Y(n7343) );
  MX4XL U10572 ( .A(\xArray[0][29] ), .B(\xArray[1][29] ), .C(\xArray[2][29] ), 
        .D(\xArray[3][29] ), .S0(n7369), .S1(n7366), .Y(n7347) );
  MX4XL U10573 ( .A(\xArray[0][30] ), .B(\xArray[1][30] ), .C(\xArray[2][30] ), 
        .D(\xArray[3][30] ), .S0(n7372), .S1(n7364), .Y(n7351) );
  MX4XL U10574 ( .A(\xArray[0][31] ), .B(\xArray[1][31] ), .C(\xArray[2][31] ), 
        .D(\xArray[3][31] ), .S0(n7373), .S1(n7365), .Y(n7355) );
  MX4XL U10575 ( .A(\xArray[4][3] ), .B(\xArray[5][3] ), .C(\xArray[6][3] ), 
        .D(\xArray[7][3] ), .S0(n7367), .S1(n7363), .Y(n7242) );
  MX4XL U10576 ( .A(\xArray[4][4] ), .B(\xArray[5][4] ), .C(\xArray[6][4] ), 
        .D(\xArray[7][4] ), .S0(n7367), .S1(n7361), .Y(n7246) );
  MX4XL U10577 ( .A(\xArray[4][5] ), .B(\xArray[5][5] ), .C(\xArray[6][5] ), 
        .D(\xArray[7][5] ), .S0(n7367), .S1(n7362), .Y(n7250) );
  MX4XL U10578 ( .A(\xArray[4][6] ), .B(\xArray[5][6] ), .C(\xArray[6][6] ), 
        .D(\xArray[7][6] ), .S0(n7368), .S1(n7362), .Y(n7254) );
  MX4XL U10579 ( .A(\xArray[4][7] ), .B(\xArray[5][7] ), .C(\xArray[6][7] ), 
        .D(\xArray[7][7] ), .S0(n7368), .S1(n7363), .Y(n7258) );
  MX4XL U10580 ( .A(\xArray[4][8] ), .B(\xArray[5][8] ), .C(\xArray[6][8] ), 
        .D(\xArray[7][8] ), .S0(n7368), .S1(n7361), .Y(n7262) );
  MX4XL U10581 ( .A(\xArray[4][9] ), .B(\xArray[5][9] ), .C(\xArray[6][9] ), 
        .D(\xArray[7][9] ), .S0(n7369), .S1(n7361), .Y(n7266) );
  MX4XL U10582 ( .A(\xArray[4][10] ), .B(\xArray[5][10] ), .C(\xArray[6][10] ), 
        .D(\xArray[7][10] ), .S0(n7369), .S1(n7361), .Y(n7270) );
  MX4XL U10583 ( .A(\xArray[4][11] ), .B(\xArray[5][11] ), .C(\xArray[6][11] ), 
        .D(\xArray[7][11] ), .S0(n7369), .S1(n7361), .Y(n7274) );
  MX4XL U10584 ( .A(\xArray[4][12] ), .B(\xArray[5][12] ), .C(\xArray[6][12] ), 
        .D(\xArray[7][12] ), .S0(n7370), .S1(n7362), .Y(n7278) );
  MX4XL U10585 ( .A(\xArray[4][13] ), .B(\xArray[5][13] ), .C(\xArray[6][13] ), 
        .D(\xArray[7][13] ), .S0(n7370), .S1(n7362), .Y(n7282) );
  MX4XL U10586 ( .A(\xArray[4][14] ), .B(\xArray[5][14] ), .C(\xArray[6][14] ), 
        .D(\xArray[7][14] ), .S0(n7370), .S1(n7362), .Y(n7286) );
  MX4XL U10587 ( .A(\xArray[4][15] ), .B(\xArray[5][15] ), .C(\xArray[6][15] ), 
        .D(\xArray[7][15] ), .S0(n7370), .S1(n7362), .Y(n7290) );
  MX4XL U10588 ( .A(\xArray[4][16] ), .B(\xArray[5][16] ), .C(\xArray[6][16] ), 
        .D(\xArray[7][16] ), .S0(n7371), .S1(n7363), .Y(n7294) );
  MX4XL U10589 ( .A(\xArray[4][17] ), .B(\xArray[5][17] ), .C(\xArray[6][17] ), 
        .D(\xArray[7][17] ), .S0(n7371), .S1(n7363), .Y(n7298) );
  MX4XL U10590 ( .A(\xArray[4][18] ), .B(\xArray[5][18] ), .C(\xArray[6][18] ), 
        .D(\xArray[7][18] ), .S0(n7371), .S1(n7363), .Y(n7302) );
  MX4XL U10591 ( .A(\xArray[4][19] ), .B(\xArray[5][19] ), .C(\xArray[6][19] ), 
        .D(\xArray[7][19] ), .S0(n7372), .S1(n7364), .Y(n7306) );
  MX4XL U10592 ( .A(\xArray[4][20] ), .B(\xArray[5][20] ), .C(\xArray[6][20] ), 
        .D(\xArray[7][20] ), .S0(n7372), .S1(n7364), .Y(n7310) );
  MX4XL U10593 ( .A(\xArray[4][21] ), .B(\xArray[5][21] ), .C(\xArray[6][21] ), 
        .D(\xArray[7][21] ), .S0(n7372), .S1(n7364), .Y(n7314) );
  MX4XL U10594 ( .A(\xArray[4][22] ), .B(\xArray[5][22] ), .C(\xArray[6][22] ), 
        .D(\xArray[7][22] ), .S0(n7373), .S1(n7365), .Y(n7318) );
  MX4XL U10595 ( .A(\xArray[4][23] ), .B(\xArray[5][23] ), .C(\xArray[6][23] ), 
        .D(\xArray[7][23] ), .S0(n7373), .S1(n7365), .Y(n7322) );
  MX4XL U10596 ( .A(\xArray[4][24] ), .B(\xArray[5][24] ), .C(\xArray[6][24] ), 
        .D(\xArray[7][24] ), .S0(n7373), .S1(n7365), .Y(n7326) );
  MX4XL U10597 ( .A(\xArray[4][25] ), .B(\xArray[5][25] ), .C(\xArray[6][25] ), 
        .D(\xArray[7][25] ), .S0(n7374), .S1(n7366), .Y(n7330) );
  MX4XL U10598 ( .A(\xArray[4][26] ), .B(\xArray[5][26] ), .C(\xArray[6][26] ), 
        .D(\xArray[7][26] ), .S0(n7374), .S1(n7366), .Y(n7334) );
  MX4XL U10599 ( .A(\xArray[4][27] ), .B(\xArray[5][27] ), .C(\xArray[6][27] ), 
        .D(\xArray[7][27] ), .S0(n7374), .S1(n7366), .Y(n7338) );
  MX4XL U10600 ( .A(\xArray[4][28] ), .B(\xArray[5][28] ), .C(\xArray[6][28] ), 
        .D(\xArray[7][28] ), .S0(n7370), .S1(n7366), .Y(n7342) );
  MX4XL U10601 ( .A(\xArray[4][29] ), .B(\xArray[5][29] ), .C(\xArray[6][29] ), 
        .D(\xArray[7][29] ), .S0(n7369), .S1(n7366), .Y(n7346) );
  MX4XL U10602 ( .A(\xArray[4][30] ), .B(\xArray[5][30] ), .C(\xArray[6][30] ), 
        .D(\xArray[7][30] ), .S0(n7372), .S1(n7364), .Y(n7350) );
  MX4XL U10603 ( .A(\xArray[4][31] ), .B(\xArray[5][31] ), .C(\xArray[6][31] ), 
        .D(\xArray[7][31] ), .S0(n7373), .S1(n7365), .Y(n7354) );
  MX4XL U10604 ( .A(\xArray[8][8] ), .B(\xArray[9][8] ), .C(\xArray[10][8] ), 
        .D(\xArray[11][8] ), .S0(n7368), .S1(n8406), .Y(n7261) );
  MX4XL U10605 ( .A(\xArray[12][8] ), .B(\xArray[13][8] ), .C(\xArray[14][8] ), 
        .D(\xArray[15][8] ), .S0(n7368), .S1(n7361), .Y(n7260) );
  MX4XL U10606 ( .A(\xArray[8][9] ), .B(\xArray[9][9] ), .C(\xArray[10][9] ), 
        .D(\xArray[11][9] ), .S0(n7369), .S1(n7361), .Y(n7265) );
  MX4XL U10607 ( .A(\xArray[12][9] ), .B(\xArray[13][9] ), .C(\xArray[14][9] ), 
        .D(\xArray[15][9] ), .S0(n7368), .S1(n7362), .Y(n7264) );
  MX4XL U10608 ( .A(\xArray[8][10] ), .B(\xArray[9][10] ), .C(\xArray[10][10] ), .D(\xArray[11][10] ), .S0(n7369), .S1(n7361), .Y(n7269) );
  MX4XL U10609 ( .A(\xArray[12][10] ), .B(\xArray[13][10] ), .C(
        \xArray[14][10] ), .D(\xArray[15][10] ), .S0(n7369), .S1(n7361), .Y(
        n7268) );
  MX4XL U10610 ( .A(\xArray[8][11] ), .B(\xArray[9][11] ), .C(\xArray[10][11] ), .D(\xArray[11][11] ), .S0(n7369), .S1(n7361), .Y(n7273) );
  MX4XL U10611 ( .A(\xArray[12][11] ), .B(\xArray[13][11] ), .C(
        \xArray[14][11] ), .D(\xArray[15][11] ), .S0(n7369), .S1(n7361), .Y(
        n7272) );
  MX4XL U10612 ( .A(\xArray[8][12] ), .B(\xArray[9][12] ), .C(\xArray[10][12] ), .D(\xArray[11][12] ), .S0(n7369), .S1(n7361), .Y(n7277) );
  MX4XL U10613 ( .A(\xArray[12][12] ), .B(\xArray[13][12] ), .C(
        \xArray[14][12] ), .D(\xArray[15][12] ), .S0(n7369), .S1(n7361), .Y(
        n7276) );
  MX4XL U10614 ( .A(\xArray[8][13] ), .B(\xArray[9][13] ), .C(\xArray[10][13] ), .D(\xArray[11][13] ), .S0(n7370), .S1(n7362), .Y(n7281) );
  MX4XL U10615 ( .A(\xArray[12][13] ), .B(\xArray[13][13] ), .C(
        \xArray[14][13] ), .D(\xArray[15][13] ), .S0(n7370), .S1(n7362), .Y(
        n7280) );
  MX4XL U10616 ( .A(\xArray[8][14] ), .B(\xArray[9][14] ), .C(\xArray[10][14] ), .D(\xArray[11][14] ), .S0(n7370), .S1(n7362), .Y(n7285) );
  MX4XL U10617 ( .A(\xArray[12][14] ), .B(\xArray[13][14] ), .C(
        \xArray[14][14] ), .D(\xArray[15][14] ), .S0(n7370), .S1(n7362), .Y(
        n7284) );
  MX4XL U10618 ( .A(\xArray[8][15] ), .B(\xArray[9][15] ), .C(\xArray[10][15] ), .D(\xArray[11][15] ), .S0(n7370), .S1(n7362), .Y(n7289) );
  MX4XL U10619 ( .A(\xArray[12][15] ), .B(\xArray[13][15] ), .C(
        \xArray[14][15] ), .D(\xArray[15][15] ), .S0(n7370), .S1(n7362), .Y(
        n7288) );
  MX4XL U10620 ( .A(\xArray[8][16] ), .B(\xArray[9][16] ), .C(\xArray[10][16] ), .D(\xArray[11][16] ), .S0(n7371), .S1(n7363), .Y(n7293) );
  MX4XL U10621 ( .A(\xArray[12][16] ), .B(\xArray[13][16] ), .C(
        \xArray[14][16] ), .D(\xArray[15][16] ), .S0(n7371), .S1(n7363), .Y(
        n7292) );
  MX4XL U10622 ( .A(\xArray[8][17] ), .B(\xArray[9][17] ), .C(\xArray[10][17] ), .D(\xArray[11][17] ), .S0(n7371), .S1(n7363), .Y(n7297) );
  MX4XL U10623 ( .A(\xArray[12][17] ), .B(\xArray[13][17] ), .C(
        \xArray[14][17] ), .D(\xArray[15][17] ), .S0(n7371), .S1(n7363), .Y(
        n7296) );
  MX4XL U10624 ( .A(\xArray[8][18] ), .B(\xArray[9][18] ), .C(\xArray[10][18] ), .D(\xArray[11][18] ), .S0(n7371), .S1(n7363), .Y(n7301) );
  MX4XL U10625 ( .A(\xArray[12][18] ), .B(\xArray[13][18] ), .C(
        \xArray[14][18] ), .D(\xArray[15][18] ), .S0(n7371), .S1(n7363), .Y(
        n7300) );
  MX4XL U10626 ( .A(\xArray[8][19] ), .B(\xArray[9][19] ), .C(\xArray[10][19] ), .D(\xArray[11][19] ), .S0(n7372), .S1(n7364), .Y(n7305) );
  MX4XL U10627 ( .A(\xArray[12][19] ), .B(\xArray[13][19] ), .C(
        \xArray[14][19] ), .D(\xArray[15][19] ), .S0(n7372), .S1(n7364), .Y(
        n7304) );
  MX4XL U10628 ( .A(\xArray[8][20] ), .B(\xArray[9][20] ), .C(\xArray[10][20] ), .D(\xArray[11][20] ), .S0(n7372), .S1(n7364), .Y(n7309) );
  MX4XL U10629 ( .A(\xArray[12][20] ), .B(\xArray[13][20] ), .C(
        \xArray[14][20] ), .D(\xArray[15][20] ), .S0(n7372), .S1(n7364), .Y(
        n7308) );
  MX4XL U10630 ( .A(\xArray[8][21] ), .B(\xArray[9][21] ), .C(\xArray[10][21] ), .D(\xArray[11][21] ), .S0(n7372), .S1(n7364), .Y(n7313) );
  MX4XL U10631 ( .A(\xArray[12][21] ), .B(\xArray[13][21] ), .C(
        \xArray[14][21] ), .D(\xArray[15][21] ), .S0(n7372), .S1(n7364), .Y(
        n7312) );
  MX4XL U10632 ( .A(\xArray[8][22] ), .B(\xArray[9][22] ), .C(\xArray[10][22] ), .D(\xArray[11][22] ), .S0(n7373), .S1(n7365), .Y(n7317) );
  MX4XL U10633 ( .A(\xArray[12][22] ), .B(\xArray[13][22] ), .C(
        \xArray[14][22] ), .D(\xArray[15][22] ), .S0(n7372), .S1(n7364), .Y(
        n7316) );
  MX4XL U10634 ( .A(\xArray[8][23] ), .B(\xArray[9][23] ), .C(\xArray[10][23] ), .D(\xArray[11][23] ), .S0(n7373), .S1(n7365), .Y(n7321) );
  MX4XL U10635 ( .A(\xArray[12][23] ), .B(\xArray[13][23] ), .C(
        \xArray[14][23] ), .D(\xArray[15][23] ), .S0(n7373), .S1(n7365), .Y(
        n7320) );
  MX4XL U10636 ( .A(\xArray[8][24] ), .B(\xArray[9][24] ), .C(\xArray[10][24] ), .D(\xArray[11][24] ), .S0(n7373), .S1(n7365), .Y(n7325) );
  MX4XL U10637 ( .A(\xArray[12][24] ), .B(\xArray[13][24] ), .C(
        \xArray[14][24] ), .D(\xArray[15][24] ), .S0(n7373), .S1(n7365), .Y(
        n7324) );
  MX4XL U10638 ( .A(\xArray[8][25] ), .B(\xArray[9][25] ), .C(\xArray[10][25] ), .D(\xArray[11][25] ), .S0(n7373), .S1(n7365), .Y(n7329) );
  MX4XL U10639 ( .A(\xArray[12][25] ), .B(\xArray[13][25] ), .C(
        \xArray[14][25] ), .D(\xArray[15][25] ), .S0(n7373), .S1(n7365), .Y(
        n7328) );
  MX4XL U10640 ( .A(\xArray[8][26] ), .B(\xArray[9][26] ), .C(\xArray[10][26] ), .D(\xArray[11][26] ), .S0(n7368), .S1(n7366), .Y(n7333) );
  MX4XL U10641 ( .A(\xArray[12][26] ), .B(\xArray[13][26] ), .C(
        \xArray[14][26] ), .D(\xArray[15][26] ), .S0(n7367), .S1(n7366), .Y(
        n7332) );
  MX4XL U10642 ( .A(\xArray[8][27] ), .B(\xArray[9][27] ), .C(\xArray[10][27] ), .D(\xArray[11][27] ), .S0(n7369), .S1(n7366), .Y(n7337) );
  MX4XL U10643 ( .A(\xArray[12][27] ), .B(\xArray[13][27] ), .C(
        \xArray[14][27] ), .D(\xArray[15][27] ), .S0(n7367), .S1(n7366), .Y(
        n7336) );
  MX4XL U10644 ( .A(\xArray[8][28] ), .B(\xArray[9][28] ), .C(\xArray[10][28] ), .D(\xArray[11][28] ), .S0(n7372), .S1(n7366), .Y(n7341) );
  MX4XL U10645 ( .A(\xArray[12][28] ), .B(\xArray[13][28] ), .C(
        \xArray[14][28] ), .D(\xArray[15][28] ), .S0(n7374), .S1(n7366), .Y(
        n7340) );
  MX4XL U10646 ( .A(\xArray[8][29] ), .B(\xArray[9][29] ), .C(\xArray[10][29] ), .D(\xArray[11][29] ), .S0(n7371), .S1(n7364), .Y(n7345) );
  MX4XL U10647 ( .A(\xArray[12][29] ), .B(\xArray[13][29] ), .C(
        \xArray[14][29] ), .D(\xArray[15][29] ), .S0(n7370), .S1(n7366), .Y(
        n7344) );
  MX4XL U10648 ( .A(\xArray[8][30] ), .B(\xArray[9][30] ), .C(\xArray[10][30] ), .D(\xArray[11][30] ), .S0(n7370), .S1(n7365), .Y(n7349) );
  MX4XL U10649 ( .A(\xArray[12][30] ), .B(\xArray[13][30] ), .C(
        \xArray[14][30] ), .D(\xArray[15][30] ), .S0(n7371), .S1(n7364), .Y(
        n7348) );
  MX4XL U10650 ( .A(\xArray[8][31] ), .B(\xArray[9][31] ), .C(\xArray[10][31] ), .D(\xArray[11][31] ), .S0(n7371), .S1(n7366), .Y(n7353) );
  MX4XL U10651 ( .A(\xArray[12][31] ), .B(\xArray[13][31] ), .C(
        \xArray[14][31] ), .D(\xArray[15][31] ), .S0(n7368), .S1(n7365), .Y(
        n7352) );
  MX4XL U10652 ( .A(\xArray[8][2] ), .B(\xArray[9][2] ), .C(\xArray[10][2] ), 
        .D(\xArray[11][2] ), .S0(outCount_next[0]), .S1(n8406), .Y(n7237) );
  MX4XL U10653 ( .A(\xArray[12][2] ), .B(\xArray[13][2] ), .C(\xArray[14][2] ), 
        .D(\xArray[15][2] ), .S0(n7367), .S1(n8406), .Y(n7236) );
  MX4XL U10654 ( .A(\xArray[8][3] ), .B(\xArray[9][3] ), .C(\xArray[10][3] ), 
        .D(\xArray[11][3] ), .S0(n7367), .S1(n8406), .Y(n7241) );
  MX4XL U10655 ( .A(\xArray[12][3] ), .B(\xArray[13][3] ), .C(\xArray[14][3] ), 
        .D(\xArray[15][3] ), .S0(n7367), .S1(n7363), .Y(n7240) );
  MX4XL U10656 ( .A(\xArray[8][4] ), .B(\xArray[9][4] ), .C(\xArray[10][4] ), 
        .D(\xArray[11][4] ), .S0(n7367), .S1(n8406), .Y(n7245) );
  MX4XL U10657 ( .A(\xArray[12][4] ), .B(\xArray[13][4] ), .C(\xArray[14][4] ), 
        .D(\xArray[15][4] ), .S0(n7367), .S1(n7361), .Y(n7244) );
  MX4XL U10658 ( .A(\xArray[8][5] ), .B(\xArray[9][5] ), .C(\xArray[10][5] ), 
        .D(\xArray[11][5] ), .S0(n7367), .S1(outCount_next[1]), .Y(n7249) );
  MX4XL U10659 ( .A(\xArray[12][5] ), .B(\xArray[13][5] ), .C(\xArray[14][5] ), 
        .D(\xArray[15][5] ), .S0(n7367), .S1(n7362), .Y(n7248) );
  MX4XL U10660 ( .A(\xArray[8][6] ), .B(\xArray[9][6] ), .C(\xArray[10][6] ), 
        .D(\xArray[11][6] ), .S0(n7368), .S1(n7361), .Y(n7253) );
  MX4XL U10661 ( .A(\xArray[12][6] ), .B(\xArray[13][6] ), .C(\xArray[14][6] ), 
        .D(\xArray[15][6] ), .S0(n7368), .S1(n7363), .Y(n7252) );
  MX4XL U10662 ( .A(\xArray[8][7] ), .B(\xArray[9][7] ), .C(\xArray[10][7] ), 
        .D(\xArray[11][7] ), .S0(n7368), .S1(n7362), .Y(n7257) );
  MX4XL U10663 ( .A(\xArray[12][7] ), .B(\xArray[13][7] ), .C(\xArray[14][7] ), 
        .D(\xArray[15][7] ), .S0(n7368), .S1(n7363), .Y(n7256) );
  MX4XL U10664 ( .A(\xArray[0][0] ), .B(\xArray[1][0] ), .C(\xArray[2][0] ), 
        .D(\xArray[3][0] ), .S0(n7374), .S1(outCount_next[1]), .Y(n7231) );
  MX4XL U10665 ( .A(\xArray[0][1] ), .B(\xArray[1][1] ), .C(\xArray[2][1] ), 
        .D(\xArray[3][1] ), .S0(n7374), .S1(n8406), .Y(n7235) );
  MX4XL U10666 ( .A(\xArray[4][0] ), .B(\xArray[5][0] ), .C(\xArray[6][0] ), 
        .D(\xArray[7][0] ), .S0(n7374), .S1(n7363), .Y(n7230) );
  MX4XL U10667 ( .A(\xArray[4][1] ), .B(\xArray[5][1] ), .C(\xArray[6][1] ), 
        .D(\xArray[7][1] ), .S0(outCount_next[0]), .S1(outCount_next[1]), .Y(
        n7234) );
  MX4XL U10668 ( .A(\xArray[4][2] ), .B(\xArray[5][2] ), .C(\xArray[6][2] ), 
        .D(\xArray[7][2] ), .S0(n7374), .S1(outCount_next[1]), .Y(n7238) );
  MX4XL U10669 ( .A(\xArray[8][0] ), .B(\xArray[9][0] ), .C(\xArray[10][0] ), 
        .D(\xArray[11][0] ), .S0(outCount_next[0]), .S1(n8406), .Y(n7229) );
  MX4XL U10670 ( .A(\xArray[12][0] ), .B(\xArray[13][0] ), .C(\xArray[14][0] ), 
        .D(\xArray[15][0] ), .S0(n7374), .S1(n8406), .Y(n7228) );
  MX4XL U10671 ( .A(\xArray[8][1] ), .B(\xArray[9][1] ), .C(\xArray[10][1] ), 
        .D(\xArray[11][1] ), .S0(n7374), .S1(n8406), .Y(n7233) );
  MX4XL U10672 ( .A(\xArray[12][1] ), .B(\xArray[13][1] ), .C(\xArray[14][1] ), 
        .D(\xArray[15][1] ), .S0(n7374), .S1(n8406), .Y(n7232) );
  AND4XL U10673 ( .A(n8407), .B(n8408), .C(n8409), .D(n8410), .Y(n8430) );
  INVXL U10674 ( .A(\xArray[4][0] ), .Y(n9393) );
  INVXL U10675 ( .A(\xArray[4][1] ), .Y(n9385) );
  INVXL U10676 ( .A(\xArray[4][2] ), .Y(n9377) );
  INVXL U10677 ( .A(\xArray[4][3] ), .Y(n9369) );
  INVXL U10678 ( .A(\xArray[4][4] ), .Y(n9361) );
  INVXL U10679 ( .A(\xArray[4][5] ), .Y(n9353) );
  INVXL U10680 ( .A(\xArray[4][6] ), .Y(n9345) );
  INVXL U10681 ( .A(\xArray[4][7] ), .Y(n9337) );
  INVXL U10682 ( .A(\xArray[4][8] ), .Y(n9329) );
  INVXL U10683 ( .A(\xArray[4][9] ), .Y(n9321) );
  INVXL U10684 ( .A(\xArray[4][10] ), .Y(n9313) );
  INVXL U10685 ( .A(\xArray[4][11] ), .Y(n9305) );
  INVXL U10686 ( .A(\xArray[4][12] ), .Y(n9297) );
  INVXL U10687 ( .A(\xArray[4][13] ), .Y(n9289) );
  INVXL U10688 ( .A(\xArray[4][14] ), .Y(n9281) );
  INVXL U10689 ( .A(\xArray[4][15] ), .Y(n9273) );
  INVXL U10690 ( .A(\xArray[4][16] ), .Y(n9265) );
  INVXL U10691 ( .A(\xArray[4][17] ), .Y(n9257) );
  INVXL U10692 ( .A(\xArray[4][18] ), .Y(n9249) );
  INVXL U10693 ( .A(\xArray[4][19] ), .Y(n9241) );
  INVXL U10694 ( .A(\xArray[4][20] ), .Y(n9233) );
  INVXL U10695 ( .A(\xArray[4][21] ), .Y(n9225) );
  INVXL U10696 ( .A(\xArray[4][22] ), .Y(n9217) );
  INVXL U10697 ( .A(\xArray[4][23] ), .Y(n9209) );
  INVXL U10698 ( .A(\xArray[4][24] ), .Y(n9201) );
  INVXL U10699 ( .A(\xArray[4][25] ), .Y(n9193) );
  INVXL U10700 ( .A(\xArray[4][26] ), .Y(n9185) );
  INVXL U10701 ( .A(\xArray[4][27] ), .Y(n9177) );
  INVXL U10702 ( .A(\xArray[4][28] ), .Y(n9169) );
  INVXL U10703 ( .A(\xArray[4][29] ), .Y(n9161) );
  INVXL U10704 ( .A(\xArray[4][30] ), .Y(n9153) );
  INVXL U10705 ( .A(\xArray[4][31] ), .Y(n9145) );
  INVXL U10706 ( .A(\xArray[15][0] ), .Y(n9391) );
  INVXL U10707 ( .A(\xArray[15][1] ), .Y(n9383) );
  INVXL U10708 ( .A(\xArray[15][2] ), .Y(n9375) );
  INVXL U10709 ( .A(\xArray[15][3] ), .Y(n9367) );
  INVXL U10710 ( .A(\xArray[15][4] ), .Y(n9359) );
  INVXL U10711 ( .A(\xArray[15][5] ), .Y(n9351) );
  INVXL U10712 ( .A(\xArray[15][6] ), .Y(n9343) );
  INVXL U10713 ( .A(\xArray[15][7] ), .Y(n9335) );
  INVXL U10714 ( .A(\xArray[15][8] ), .Y(n9327) );
  INVXL U10715 ( .A(\xArray[15][9] ), .Y(n9319) );
  INVXL U10716 ( .A(\xArray[15][10] ), .Y(n9311) );
  INVXL U10717 ( .A(\xArray[15][11] ), .Y(n9303) );
  INVXL U10718 ( .A(\xArray[15][12] ), .Y(n9295) );
  INVXL U10719 ( .A(\xArray[15][13] ), .Y(n9287) );
  INVXL U10720 ( .A(\xArray[15][14] ), .Y(n9279) );
  INVXL U10721 ( .A(\xArray[15][15] ), .Y(n9271) );
  INVXL U10722 ( .A(\xArray[15][16] ), .Y(n9263) );
  INVXL U10723 ( .A(\xArray[15][17] ), .Y(n9255) );
  INVXL U10724 ( .A(\xArray[15][18] ), .Y(n9247) );
  INVXL U10725 ( .A(\xArray[15][19] ), .Y(n9239) );
  INVXL U10726 ( .A(\xArray[15][20] ), .Y(n9231) );
  INVXL U10727 ( .A(\xArray[15][21] ), .Y(n9223) );
  INVXL U10728 ( .A(\xArray[15][22] ), .Y(n9215) );
  INVXL U10729 ( .A(\xArray[15][23] ), .Y(n9207) );
  INVXL U10730 ( .A(\xArray[15][24] ), .Y(n9199) );
  INVXL U10731 ( .A(\xArray[15][25] ), .Y(n9191) );
  INVXL U10732 ( .A(\xArray[15][26] ), .Y(n9183) );
  INVXL U10733 ( .A(\xArray[15][27] ), .Y(n9175) );
  INVXL U10734 ( .A(\xArray[15][28] ), .Y(n9167) );
  INVXL U10735 ( .A(\xArray[15][29] ), .Y(n9159) );
  INVXL U10736 ( .A(\xArray[15][30] ), .Y(n9151) );
  INVXL U10737 ( .A(\xArray[15][31] ), .Y(n9143) );
  INVXL U10738 ( .A(\xArray[4][32] ), .Y(n9137) );
  INVXL U10739 ( .A(\xArray[4][33] ), .Y(n9129) );
  INVXL U10740 ( .A(\xArray[4][34] ), .Y(n9121) );
  INVXL U10741 ( .A(\xArray[4][35] ), .Y(n9113) );
  INVXL U10742 ( .A(\xArray[4][36] ), .Y(n9105) );
  INVXL U10743 ( .A(\xArray[4][37] ), .Y(n9097) );
  INVXL U10744 ( .A(\xArray[4][38] ), .Y(n9089) );
  INVXL U10745 ( .A(\xArray[4][39] ), .Y(n9081) );
  INVXL U10746 ( .A(\xArray[4][40] ), .Y(n9073) );
  INVXL U10747 ( .A(\xArray[4][41] ), .Y(n9065) );
  INVXL U10748 ( .A(\xArray[15][32] ), .Y(n9135) );
  INVXL U10749 ( .A(\xArray[15][33] ), .Y(n9127) );
  INVXL U10750 ( .A(\xArray[15][34] ), .Y(n9119) );
  INVXL U10751 ( .A(\xArray[15][35] ), .Y(n9111) );
  INVXL U10752 ( .A(\xArray[15][36] ), .Y(n9103) );
  INVXL U10753 ( .A(\xArray[15][37] ), .Y(n9095) );
  INVXL U10754 ( .A(\xArray[15][38] ), .Y(n9087) );
  INVXL U10755 ( .A(\xArray[15][39] ), .Y(n9079) );
  INVXL U10756 ( .A(\xArray[15][40] ), .Y(n9071) );
  INVXL U10757 ( .A(\xArray[15][41] ), .Y(n9063) );
  INVX3 U10758 ( .A(b_in[0]), .Y(n8845) );
  INVX3 U10759 ( .A(b_in[1]), .Y(n8844) );
  INVX3 U10760 ( .A(b_in[2]), .Y(n8843) );
  INVX3 U10761 ( .A(b_in[3]), .Y(n8842) );
  INVX3 U10762 ( .A(b_in[4]), .Y(n8841) );
  INVX3 U10763 ( .A(b_in[5]), .Y(n8840) );
  INVX3 U10764 ( .A(b_in[6]), .Y(n8839) );
  INVX3 U10765 ( .A(b_in[7]), .Y(n8838) );
  INVX3 U10766 ( .A(b_in[8]), .Y(n8837) );
  INVX3 U10767 ( .A(b_in[9]), .Y(n8836) );
  INVX3 U10768 ( .A(b_in[10]), .Y(n8835) );
  INVX3 U10769 ( .A(b_in[11]), .Y(n8834) );
  INVX3 U10770 ( .A(b_in[12]), .Y(n8833) );
  INVX3 U10771 ( .A(b_in[13]), .Y(n8832) );
  INVX3 U10772 ( .A(b_in[14]), .Y(n8831) );
  CLKINVX1 U10773 ( .A(reset), .Y(n8830) );
  OR2X1 U10774 ( .A(n8315), .B(n1544), .Y(n6715) );
  OR2X1 U10775 ( .A(n7719), .B(n1546), .Y(n6716) );
  NAND3X6 U10776 ( .A(n6715), .B(n6716), .C(n1738), .Y(N33771) );
  OA22X4 U10777 ( .A0(n7756), .A1(n1287), .B0(n8345), .B1(n1739), .Y(n1738) );
  CLKBUFX3 U10778 ( .A(n6589), .Y(n8012) );
  CLKBUFX3 U10779 ( .A(n6577), .Y(n8025) );
  CLKBUFX3 U10780 ( .A(n6578), .Y(n8089) );
  CLKBUFX3 U10781 ( .A(n6589), .Y(n8011) );
  CLKBUFX3 U10782 ( .A(n6577), .Y(n8024) );
  CLKBUFX3 U10783 ( .A(n6590), .Y(n8076) );
  CLKBUFX3 U10784 ( .A(n6578), .Y(n8088) );
  CLKBUFX3 U10785 ( .A(n6590), .Y(n8075) );
  CLKBUFX3 U10786 ( .A(n6589), .Y(n8010) );
  CLKBUFX3 U10787 ( .A(n6577), .Y(n8023) );
  CLKBUFX3 U10788 ( .A(n6590), .Y(n8074) );
  CLKBUFX3 U10789 ( .A(n6578), .Y(n8087) );
  CLKBUFX3 U10790 ( .A(n6580), .Y(n8166) );
  CLKBUFX3 U10791 ( .A(n8164), .Y(n8165) );
  CLKBUFX3 U10792 ( .A(n6581), .Y(n8000) );
  CLKBUFX3 U10793 ( .A(n6575), .Y(n8038) );
  CLKBUFX3 U10794 ( .A(n6587), .Y(n8153) );
  CLKBUFX3 U10795 ( .A(n6581), .Y(n7999) );
  CLKBUFX3 U10796 ( .A(n6575), .Y(n8037) );
  CLKBUFX3 U10797 ( .A(n6587), .Y(n8152) );
  CLKBUFX3 U10798 ( .A(n6581), .Y(n7998) );
  CLKBUFX3 U10799 ( .A(n6575), .Y(n8036) );
  CLKBUFX3 U10800 ( .A(n6587), .Y(n8151) );
  INVX3 U10801 ( .A(n7779), .Y(n7768) );
  INVX4 U10802 ( .A(n7775), .Y(n7772) );
  INVX4 U10803 ( .A(n7776), .Y(n7771) );
  INVX3 U10804 ( .A(n7774), .Y(n7773) );
  INVX3 U10805 ( .A(n7778), .Y(n7769) );
  INVX3 U10806 ( .A(n7778), .Y(n7770) );
  INVX3 U10807 ( .A(n7816), .Y(n7809) );
  INVX3 U10808 ( .A(n7915), .Y(n7911) );
  INVX3 U10809 ( .A(n7897), .Y(n7891) );
  INVX3 U10810 ( .A(n7820), .Y(n7808) );
  INVX3 U10811 ( .A(n7915), .Y(n7910) );
  INVX3 U10812 ( .A(n7916), .Y(n7909) );
  INVX3 U10813 ( .A(n7901), .Y(n7890) );
  CLKINVX1 U10814 ( .A(n7496), .Y(n8453) );
  CLKINVX1 U10815 ( .A(n7500), .Y(n8458) );
  CLKINVX1 U10816 ( .A(n7498), .Y(n8448) );
  INVX3 U10817 ( .A(n6693), .Y(n8187) );
  INVX3 U10818 ( .A(n8205), .Y(n8189) );
  INVX3 U10819 ( .A(n8202), .Y(n8196) );
  INVX3 U10820 ( .A(n8206), .Y(n8186) );
  INVX3 U10821 ( .A(n8205), .Y(n8190) );
  INVX3 U10822 ( .A(n8204), .Y(n8192) );
  AO22X1 U10823 ( .A0(N29671), .A1(n7773), .B0(N30439), .B1(n7793), .Y(n3738)
         );
  AO22X1 U10824 ( .A0(N29672), .A1(n7773), .B0(N30440), .B1(n7793), .Y(n3720)
         );
  AO22X1 U10825 ( .A0(N29673), .A1(n7773), .B0(N30441), .B1(n7790), .Y(n3699)
         );
  AO22X1 U10826 ( .A0(N29666), .A1(n7773), .B0(N30434), .B1(n7793), .Y(n3828)
         );
  AO22X1 U10827 ( .A0(N29665), .A1(n7772), .B0(N30433), .B1(n7793), .Y(n3846)
         );
  AO22X1 U10828 ( .A0(N29668), .A1(n7772), .B0(N30436), .B1(n7793), .Y(n3792)
         );
  INVX3 U10829 ( .A(n8207), .Y(n8184) );
  AO22X1 U10830 ( .A0(N29662), .A1(n7772), .B0(N30430), .B1(n7793), .Y(n3900)
         );
  AO22X1 U10831 ( .A0(N29663), .A1(n7772), .B0(N30431), .B1(n7793), .Y(n3882)
         );
  AO22X1 U10832 ( .A0(N29660), .A1(n7771), .B0(N30428), .B1(n7793), .Y(n3936)
         );
  CLKBUFX3 U10833 ( .A(n1747), .Y(n8176) );
  CLKBUFX3 U10834 ( .A(n1746), .Y(n8180) );
  AO22X1 U10835 ( .A0(N29657), .A1(n7771), .B0(N30425), .B1(n7793), .Y(n3990)
         );
  AO22X1 U10836 ( .A0(N29658), .A1(n7771), .B0(N30426), .B1(n7793), .Y(n3972)
         );
  INVX3 U10837 ( .A(n8276), .Y(n8253) );
  INVX3 U10838 ( .A(n8205), .Y(n8188) );
  AO22X1 U10839 ( .A0(N29654), .A1(n7772), .B0(N30422), .B1(n7792), .Y(n4044)
         );
  AO22X1 U10840 ( .A0(N29655), .A1(n7771), .B0(N30423), .B1(n7792), .Y(n4026)
         );
  INVX3 U10841 ( .A(n8203), .Y(n8195) );
  INVX3 U10842 ( .A(n8204), .Y(n8191) );
  AO22X1 U10843 ( .A0(N29651), .A1(n7771), .B0(N30419), .B1(n7792), .Y(n4098)
         );
  AO22X1 U10844 ( .A0(N29652), .A1(n7771), .B0(N30420), .B1(n7792), .Y(n4080)
         );
  AO22X1 U10845 ( .A0(N29647), .A1(n7771), .B0(N30415), .B1(n7792), .Y(n4170)
         );
  AO22X1 U10846 ( .A0(N29649), .A1(n7771), .B0(N30417), .B1(n7792), .Y(n4134)
         );
  AO22X1 U10847 ( .A0(N29650), .A1(n7771), .B0(N30418), .B1(n7792), .Y(n4116)
         );
  INVX3 U10848 ( .A(n8202), .Y(n8197) );
  AO22X1 U10849 ( .A0(N29644), .A1(n7771), .B0(N30412), .B1(n7792), .Y(n4224)
         );
  AO22X1 U10850 ( .A0(N29646), .A1(n7771), .B0(N30414), .B1(n7792), .Y(n4188)
         );
  AO22X1 U10851 ( .A0(N29641), .A1(n7771), .B0(N30409), .B1(n7792), .Y(n4278)
         );
  AO22X1 U10852 ( .A0(N29642), .A1(n7771), .B0(N30410), .B1(n7792), .Y(n4260)
         );
  AO22X1 U10853 ( .A0(N29639), .A1(n7771), .B0(N30407), .B1(n7792), .Y(n4314)
         );
  AO22X1 U10854 ( .A0(N29636), .A1(n7771), .B0(N30404), .B1(n7791), .Y(n4368)
         );
  AO22X1 U10855 ( .A0(N29637), .A1(n7771), .B0(N30405), .B1(n7791), .Y(n4350)
         );
  AO22X1 U10856 ( .A0(N29634), .A1(n7772), .B0(N30402), .B1(n7791), .Y(n4404)
         );
  AO22X1 U10857 ( .A0(N29631), .A1(n7772), .B0(N30399), .B1(n7791), .Y(n4458)
         );
  AO22X1 U10858 ( .A0(N29633), .A1(n7771), .B0(N30401), .B1(n7791), .Y(n4422)
         );
  INVX3 U10859 ( .A(n8206), .Y(n8185) );
  AO22X1 U10860 ( .A0(N29628), .A1(n7772), .B0(N30396), .B1(n7791), .Y(n4512)
         );
  AO22X1 U10861 ( .A0(N29629), .A1(n7772), .B0(N30397), .B1(n7791), .Y(n4494)
         );
  CLKBUFX3 U10862 ( .A(n1746), .Y(n8179) );
  AO22X1 U10863 ( .A0(N29624), .A1(n7772), .B0(N30392), .B1(n7791), .Y(n4584)
         );
  AO22X1 U10864 ( .A0(N29626), .A1(n7772), .B0(N30394), .B1(n7790), .Y(n4548)
         );
  AO22X1 U10865 ( .A0(N29622), .A1(n7772), .B0(N30390), .B1(n7791), .Y(n4620)
         );
  AO22X1 U10866 ( .A0(N29617), .A1(n7773), .B0(N30385), .B1(n7790), .Y(n4710)
         );
  AO22X1 U10867 ( .A0(N29620), .A1(n7773), .B0(N30388), .B1(n7790), .Y(n4656)
         );
  AO22X1 U10868 ( .A0(N29621), .A1(n7772), .B0(N30389), .B1(n7791), .Y(n4638)
         );
  AO22X1 U10869 ( .A0(N29618), .A1(n7773), .B0(N30386), .B1(n7791), .Y(n4692)
         );
  AO22X1 U10870 ( .A0(N29619), .A1(n7773), .B0(N30387), .B1(n7790), .Y(n4674)
         );
  AO22X1 U10871 ( .A0(N29615), .A1(n7773), .B0(N30383), .B1(n7791), .Y(n4746)
         );
  AO22X1 U10872 ( .A0(N29614), .A1(n7773), .B0(N30382), .B1(n7790), .Y(n4764)
         );
  AO22X1 U10873 ( .A0(N29611), .A1(n7773), .B0(N30379), .B1(n7790), .Y(n4818)
         );
  AO22X1 U10874 ( .A0(N29612), .A1(n7773), .B0(N30380), .B1(n7790), .Y(n4800)
         );
  AO22X1 U10875 ( .A0(N29613), .A1(n7773), .B0(N30381), .B1(n7790), .Y(n4782)
         );
  INVX3 U10876 ( .A(n8204), .Y(n8193) );
  INVX3 U10877 ( .A(n8203), .Y(n8194) );
  CLKBUFX3 U10878 ( .A(n8173), .Y(n8174) );
  CLKBUFX3 U10879 ( .A(n7981), .Y(n7984) );
  CLKBUFX3 U10880 ( .A(n7981), .Y(n7983) );
  CLKBUFX3 U10881 ( .A(n8109), .Y(n8112) );
  CLKBUFX3 U10882 ( .A(n7981), .Y(n7982) );
  CLKBUFX3 U10883 ( .A(n8109), .Y(n8111) );
  CLKBUFX3 U10884 ( .A(n8058), .Y(n8060) );
  CLKBUFX3 U10885 ( .A(n2599), .Y(n8137) );
  CLKBUFX3 U10886 ( .A(n8058), .Y(n8059) );
  CLKBUFX3 U10887 ( .A(n2599), .Y(n8136) );
  CLKBUFX3 U10888 ( .A(n2599), .Y(n8135) );
  CLKBUFX3 U10889 ( .A(n3572), .Y(n7980) );
  CLKBUFX3 U10890 ( .A(n2808), .Y(n8108) );
  CLKBUFX3 U10891 ( .A(n3572), .Y(n7979) );
  CLKBUFX3 U10892 ( .A(n2808), .Y(n8107) );
  CLKBUFX3 U10893 ( .A(n3572), .Y(n7978) );
  CLKBUFX3 U10894 ( .A(n2808), .Y(n8106) );
  AND2X2 U10895 ( .A(n7986), .B(n7989), .Y(n3636) );
  AND2X2 U10896 ( .A(n8050), .B(n8053), .Y(n3290) );
  AND2X2 U10897 ( .A(n8101), .B(n8104), .Y(n3007) );
  AND2X2 U10898 ( .A(n8114), .B(n8117), .Y(n2935) );
  AND2X2 U10899 ( .A(n8127), .B(n8129), .Y(n2800) );
  AND2X2 U10900 ( .A(n8062), .B(n8064), .Y(n3218) );
  AND2X2 U10901 ( .A(n8139), .B(n8141), .Y(n2728) );
  CLKBUFX3 U10902 ( .A(n6580), .Y(n8164) );
  INVX3 U10903 ( .A(n7881), .Y(n7868) );
  CLKBUFX3 U10904 ( .A(n7780), .Y(n7779) );
  CLKBUFX3 U10905 ( .A(n3671), .Y(n7937) );
  CLKBUFX3 U10906 ( .A(n7935), .Y(n7936) );
  CLKBUFX3 U10907 ( .A(n6604), .Y(n7940) );
  CLKBUFX3 U10908 ( .A(n6604), .Y(n7939) );
  CLKBUFX3 U10909 ( .A(n6604), .Y(n7938) );
  INVX3 U10910 ( .A(n7879), .Y(n7872) );
  INVX3 U10911 ( .A(n7878), .Y(n7873) );
  INVX3 U10912 ( .A(n7877), .Y(n7874) );
  CLKBUFX3 U10913 ( .A(n7781), .Y(n7776) );
  CLKBUFX3 U10914 ( .A(n7782), .Y(n7775) );
  CLKBUFX3 U10915 ( .A(n7782), .Y(n7774) );
  INVX3 U10916 ( .A(n7797), .Y(n7790) );
  CLKBUFX3 U10917 ( .A(n3498), .Y(n8004) );
  CLKBUFX3 U10918 ( .A(n8006), .Y(n8005) );
  CLKBUFX3 U10919 ( .A(n3660), .Y(n7961) );
  CLKBUFX3 U10920 ( .A(n3660), .Y(n7960) );
  CLKBUFX3 U10921 ( .A(n3660), .Y(n7959) );
  INVX3 U10922 ( .A(n7794), .Y(n7793) );
  CLKBUFX3 U10923 ( .A(n7944), .Y(n7946) );
  CLKBUFX3 U10924 ( .A(n7944), .Y(n7945) );
  CLKBUFX3 U10925 ( .A(n7962), .Y(n7965) );
  CLKBUFX3 U10926 ( .A(n7962), .Y(n7964) );
  CLKBUFX3 U10927 ( .A(n7962), .Y(n7963) );
  CLKBUFX3 U10928 ( .A(n3663), .Y(n7954) );
  CLKBUFX3 U10929 ( .A(n3663), .Y(n7953) );
  CLKINVX1 U10930 ( .A(n7876), .Y(n7875) );
  CLKBUFX3 U10931 ( .A(n3663), .Y(n7955) );
  INVX3 U10932 ( .A(n7880), .Y(n7869) );
  INVX3 U10933 ( .A(n7880), .Y(n7870) );
  INVX3 U10934 ( .A(n7882), .Y(n7871) );
  CLKBUFX3 U10935 ( .A(n7928), .Y(n7915) );
  CLKBUFX3 U10936 ( .A(n7826), .Y(n7814) );
  CLKBUFX3 U10937 ( .A(n7928), .Y(n7916) );
  CLKBUFX3 U10938 ( .A(n7780), .Y(n7778) );
  CLKBUFX3 U10939 ( .A(n7781), .Y(n7777) );
  INVX3 U10940 ( .A(n7813), .Y(n7811) );
  INVX3 U10941 ( .A(n7928), .Y(n7913) );
  INVX3 U10942 ( .A(n7897), .Y(n7893) );
  INVX3 U10943 ( .A(n7815), .Y(n7810) );
  INVX3 U10944 ( .A(n7928), .Y(n7912) );
  INVX3 U10945 ( .A(n7908), .Y(n7892) );
  INVX3 U10946 ( .A(n7802), .Y(n7789) );
  INVX3 U10947 ( .A(n7835), .Y(n7829) );
  INVX3 U10948 ( .A(n7854), .Y(n7848) );
  INVX3 U10949 ( .A(n7801), .Y(n7788) );
  INVX3 U10950 ( .A(n7802), .Y(n7787) );
  INVX3 U10951 ( .A(n7836), .Y(n7828) );
  INVX3 U10952 ( .A(n7801), .Y(n7786) );
  INVX3 U10953 ( .A(n7802), .Y(n7785) );
  CLKBUFX3 U10954 ( .A(n7825), .Y(n7815) );
  CLKBUFX3 U10955 ( .A(n7902), .Y(n7895) );
  CLKBUFX3 U10956 ( .A(n7825), .Y(n7816) );
  CLKBUFX3 U10957 ( .A(n7902), .Y(n7896) );
  CLKBUFX3 U10958 ( .A(n7825), .Y(n7817) );
  CLKBUFX3 U10959 ( .A(n7928), .Y(n7917) );
  CLKBUFX3 U10960 ( .A(n7889), .Y(n7897) );
  CLKBUFX3 U10961 ( .A(n7826), .Y(n7818) );
  CLKBUFX3 U10962 ( .A(n7928), .Y(n7918) );
  CLKBUFX3 U10963 ( .A(n7908), .Y(n7898) );
  CLKBUFX3 U10964 ( .A(n7927), .Y(n7919) );
  CLKBUFX3 U10965 ( .A(n7908), .Y(n7899) );
  CLKBUFX3 U10966 ( .A(n7824), .Y(n7819) );
  CLKBUFX3 U10967 ( .A(n7927), .Y(n7920) );
  CLKBUFX3 U10968 ( .A(n7908), .Y(n7900) );
  CLKBUFX3 U10969 ( .A(n7824), .Y(n7820) );
  CLKBUFX3 U10970 ( .A(n7927), .Y(n7921) );
  CLKBUFX3 U10971 ( .A(n7897), .Y(n7901) );
  CLKBUFX3 U10972 ( .A(n7927), .Y(n7922) );
  CLKBUFX3 U10973 ( .A(n7889), .Y(n7902) );
  CLKBUFX3 U10974 ( .A(n7901), .Y(n7903) );
  CLKBUFX3 U10975 ( .A(n7906), .Y(n7904) );
  CLKBUFX3 U10976 ( .A(n7926), .Y(n7923) );
  CLKBUFX3 U10977 ( .A(n7907), .Y(n7905) );
  CLKBUFX3 U10978 ( .A(n7823), .Y(n7821) );
  CLKBUFX3 U10979 ( .A(n7926), .Y(n7924) );
  CLKBUFX3 U10980 ( .A(n7908), .Y(n7906) );
  CLKBUFX3 U10981 ( .A(n7823), .Y(n7822) );
  CLKBUFX3 U10982 ( .A(n7926), .Y(n7925) );
  CLKBUFX3 U10983 ( .A(n7908), .Y(n7907) );
  CLKINVX1 U10984 ( .A(n7823), .Y(n7812) );
  CLKINVX1 U10985 ( .A(n3678), .Y(n7914) );
  CLKINVX1 U10986 ( .A(n7902), .Y(n7894) );
  NAND2X1 U10987 ( .A(n3736), .B(n3737), .Y(n2605) );
  AOI222XL U10988 ( .A0(N34791), .A1(n7765), .B0(N32743), .B1(n7706), .C0(
        N31975), .C1(n7763), .Y(n3736) );
  CLKBUFX3 U10989 ( .A(n2607), .Y(n7494) );
  NAND2X1 U10990 ( .A(n3754), .B(n3755), .Y(n2607) );
  AOI222XL U10991 ( .A0(N34790), .A1(n7764), .B0(N32742), .B1(n7706), .C0(
        N31974), .C1(n7763), .Y(n3754) );
  AOI221XL U10992 ( .A0(N33702), .A1(n7874), .B0(N31398), .B1(n7703), .C0(
        n3756), .Y(n3755) );
  NAND2X1 U10993 ( .A(n3696), .B(n3697), .Y(n2600) );
  AOI222XL U10994 ( .A0(N34793), .A1(n7764), .B0(N32745), .B1(n7704), .C0(
        N31977), .C1(n7761), .Y(n3696) );
  CLKBUFX3 U10995 ( .A(n2615), .Y(n7486) );
  NAND2X1 U10996 ( .A(n3826), .B(n3827), .Y(n2615) );
  AOI222XL U10997 ( .A0(N34786), .A1(n7766), .B0(N32738), .B1(n7706), .C0(
        N31970), .C1(n7763), .Y(n3826) );
  AOI221XL U10998 ( .A0(N33698), .A1(n7874), .B0(N31394), .B1(n7702), .C0(
        n3828), .Y(n3827) );
  CLKBUFX3 U10999 ( .A(n2613), .Y(n7488) );
  NAND2X1 U11000 ( .A(n3808), .B(n3809), .Y(n2613) );
  AOI222XL U11001 ( .A0(N34787), .A1(n7765), .B0(N32739), .B1(n7706), .C0(
        N31971), .C1(n7763), .Y(n3808) );
  AOI221XL U11002 ( .A0(N33699), .A1(n7874), .B0(N31395), .B1(n7702), .C0(
        n3810), .Y(n3809) );
  CLKBUFX3 U11003 ( .A(n2611), .Y(n7490) );
  NAND2X1 U11004 ( .A(n3790), .B(n3791), .Y(n2611) );
  AOI222XL U11005 ( .A0(N34788), .A1(n7765), .B0(N32740), .B1(n7706), .C0(
        N31972), .C1(n7763), .Y(n3790) );
  AOI221XL U11006 ( .A0(N33700), .A1(n7874), .B0(N31396), .B1(n7703), .C0(
        n3792), .Y(n3791) );
  CLKBUFX3 U11007 ( .A(n2609), .Y(n7492) );
  NAND2X1 U11008 ( .A(n3772), .B(n3773), .Y(n2609) );
  AOI222XL U11009 ( .A0(N34789), .A1(n3700), .B0(N32741), .B1(n7706), .C0(
        N31973), .C1(n7763), .Y(n3772) );
  AOI221XL U11010 ( .A0(N33701), .A1(n7874), .B0(N31397), .B1(n7703), .C0(
        n3774), .Y(n3773) );
  NAND2X1 U11011 ( .A(n3718), .B(n3719), .Y(n2603) );
  AOI222XL U11012 ( .A0(N34792), .A1(n7764), .B0(N32744), .B1(n7706), .C0(
        N31976), .C1(n7763), .Y(n3718) );
  CLKBUFX3 U11013 ( .A(n7745), .Y(n7758) );
  CLKBUFX3 U11014 ( .A(n7747), .Y(n7760) );
  INVX3 U11015 ( .A(n8275), .Y(n8268) );
  INVX3 U11016 ( .A(n8275), .Y(n8270) );
  INVX3 U11017 ( .A(n8274), .Y(n8273) );
  CLKBUFX3 U11018 ( .A(n7735), .Y(n7723) );
  CLKBUFX3 U11019 ( .A(n2623), .Y(n7478) );
  NAND2X1 U11020 ( .A(n3898), .B(n3899), .Y(n2623) );
  AOI222XL U11021 ( .A0(N34782), .A1(n7766), .B0(N32734), .B1(n7706), .C0(
        N31966), .C1(n7763), .Y(n3898) );
  AOI221XL U11022 ( .A0(N33694), .A1(n7873), .B0(N31390), .B1(n7702), .C0(
        n3900), .Y(n3899) );
  CLKBUFX3 U11023 ( .A(n2621), .Y(n7480) );
  NAND2X1 U11024 ( .A(n3880), .B(n3881), .Y(n2621) );
  AOI222XL U11025 ( .A0(N34783), .A1(n7765), .B0(N32735), .B1(n7706), .C0(
        N31967), .C1(n7763), .Y(n3880) );
  AOI221XL U11026 ( .A0(N33695), .A1(n7873), .B0(N31391), .B1(n7702), .C0(
        n3882), .Y(n3881) );
  CLKBUFX3 U11027 ( .A(n2619), .Y(n7482) );
  NAND2X1 U11028 ( .A(n3862), .B(n3863), .Y(n2619) );
  AOI222XL U11029 ( .A0(N34784), .A1(n7766), .B0(N32736), .B1(n7706), .C0(
        N31968), .C1(n7763), .Y(n3862) );
  AOI221XL U11030 ( .A0(N33696), .A1(n7874), .B0(N31392), .B1(n7702), .C0(
        n3864), .Y(n3863) );
  CLKBUFX3 U11031 ( .A(n2617), .Y(n7484) );
  NAND2X1 U11032 ( .A(n3844), .B(n3845), .Y(n2617) );
  AOI222XL U11033 ( .A0(N34785), .A1(n7765), .B0(N32737), .B1(n7706), .C0(
        N31969), .C1(n7763), .Y(n3844) );
  AOI221XL U11034 ( .A0(N33697), .A1(n7873), .B0(N31393), .B1(n7702), .C0(
        n3846), .Y(n3845) );
  CLKBUFX3 U11035 ( .A(n7743), .Y(n7753) );
  CLKBUFX3 U11036 ( .A(n7743), .Y(n7754) );
  CLKBUFX3 U11037 ( .A(n7749), .Y(n7756) );
  INVX3 U11038 ( .A(n8274), .Y(n8272) );
  CLKBUFX3 U11039 ( .A(n7734), .Y(n7724) );
  CLKBUFX3 U11040 ( .A(n7738), .Y(n7716) );
  INVX3 U11041 ( .A(n8326), .Y(n8315) );
  CLKBUFX3 U11042 ( .A(n2625), .Y(n7476) );
  NAND2X1 U11043 ( .A(n3916), .B(n3917), .Y(n2625) );
  AOI222XL U11044 ( .A0(N34781), .A1(n7765), .B0(N32733), .B1(n7706), .C0(
        N31965), .C1(n7763), .Y(n3916) );
  AOI221XL U11045 ( .A0(N33693), .A1(n7873), .B0(N31389), .B1(n7702), .C0(
        n3918), .Y(n3917) );
  CLKBUFX3 U11046 ( .A(n2629), .Y(n7472) );
  NAND2X1 U11047 ( .A(n3952), .B(n3953), .Y(n2629) );
  AOI222XL U11048 ( .A0(N34779), .A1(n7766), .B0(N32731), .B1(n7706), .C0(
        N31963), .C1(n7762), .Y(n3952) );
  AOI221XL U11049 ( .A0(N33691), .A1(n7873), .B0(N31387), .B1(n7702), .C0(
        n3954), .Y(n3953) );
  CLKBUFX3 U11050 ( .A(n2627), .Y(n7474) );
  NAND2X1 U11051 ( .A(n3934), .B(n3935), .Y(n2627) );
  AOI222XL U11052 ( .A0(N34780), .A1(n3700), .B0(N32732), .B1(n7706), .C0(
        N31964), .C1(n7763), .Y(n3934) );
  AOI221XL U11053 ( .A0(N33692), .A1(n7872), .B0(N31388), .B1(n7702), .C0(
        n3936), .Y(n3935) );
  CLKBUFX3 U11054 ( .A(n2639), .Y(n7462) );
  NAND2X1 U11055 ( .A(n4042), .B(n4043), .Y(n2639) );
  AOI222XL U11056 ( .A0(N34774), .A1(n7764), .B0(N32726), .B1(n7705), .C0(
        N31958), .C1(n7762), .Y(n4042) );
  AOI221XL U11057 ( .A0(N33686), .A1(n7873), .B0(N31382), .B1(n7702), .C0(
        n4044), .Y(n4043) );
  CLKBUFX3 U11058 ( .A(n2637), .Y(n7464) );
  NAND2X1 U11059 ( .A(n4024), .B(n4025), .Y(n2637) );
  AOI222XL U11060 ( .A0(N34775), .A1(n7764), .B0(N32727), .B1(n7706), .C0(
        N31959), .C1(n7762), .Y(n4024) );
  AOI221XL U11061 ( .A0(N33687), .A1(n7872), .B0(N31383), .B1(n7702), .C0(
        n4026), .Y(n4025) );
  CLKBUFX3 U11062 ( .A(n2635), .Y(n7466) );
  NAND2X1 U11063 ( .A(n4006), .B(n4007), .Y(n2635) );
  AOI222XL U11064 ( .A0(N34776), .A1(n7765), .B0(N32728), .B1(n7706), .C0(
        N31960), .C1(n7762), .Y(n4006) );
  AOI221XL U11065 ( .A0(N33688), .A1(n7873), .B0(N31384), .B1(n7702), .C0(
        n4008), .Y(n4007) );
  CLKBUFX3 U11066 ( .A(n2633), .Y(n7468) );
  NAND2X1 U11067 ( .A(n3988), .B(n3989), .Y(n2633) );
  AOI222XL U11068 ( .A0(N34777), .A1(n7766), .B0(N32729), .B1(n7706), .C0(
        N31961), .C1(n7762), .Y(n3988) );
  AOI221XL U11069 ( .A0(N33689), .A1(n7872), .B0(N31385), .B1(n7702), .C0(
        n3990), .Y(n3989) );
  CLKBUFX3 U11070 ( .A(n2631), .Y(n7470) );
  NAND2X1 U11071 ( .A(n3970), .B(n3971), .Y(n2631) );
  AOI222XL U11072 ( .A0(N34778), .A1(n7764), .B0(N32730), .B1(n7706), .C0(
        N31962), .C1(n7762), .Y(n3970) );
  AOI221XL U11073 ( .A0(N33690), .A1(n7873), .B0(N31386), .B1(n7702), .C0(
        n3972), .Y(n3971) );
  CLKBUFX3 U11074 ( .A(n7744), .Y(n7755) );
  CLKBUFX3 U11075 ( .A(n7745), .Y(n7757) );
  CLKBUFX3 U11076 ( .A(n7746), .Y(n7759) );
  CLKBUFX3 U11077 ( .A(n8217), .Y(n8208) );
  CLKBUFX3 U11078 ( .A(n2645), .Y(n7457) );
  NAND2X1 U11079 ( .A(n4096), .B(n4097), .Y(n2645) );
  AOI222XL U11080 ( .A0(N34771), .A1(n7766), .B0(N32723), .B1(n8857), .C0(
        N31955), .C1(n7762), .Y(n4096) );
  AOI221XL U11081 ( .A0(N33683), .A1(n7872), .B0(N31379), .B1(n7702), .C0(
        n4098), .Y(n4097) );
  CLKBUFX3 U11082 ( .A(n2643), .Y(n7459) );
  NAND2X1 U11083 ( .A(n4078), .B(n4079), .Y(n2643) );
  AOI222XL U11084 ( .A0(N34772), .A1(n7764), .B0(N32724), .B1(n8857), .C0(
        N31956), .C1(n7762), .Y(n4078) );
  AOI221XL U11085 ( .A0(N33684), .A1(n7872), .B0(N31380), .B1(n7702), .C0(
        n4080), .Y(n4079) );
  CLKBUFX3 U11086 ( .A(n2641), .Y(n7461) );
  NAND2X1 U11087 ( .A(n4060), .B(n4061), .Y(n2641) );
  AOI222XL U11088 ( .A0(N34773), .A1(n3700), .B0(N32725), .B1(n8857), .C0(
        N31957), .C1(n7762), .Y(n4060) );
  AOI221XL U11089 ( .A0(N33685), .A1(n7872), .B0(N31381), .B1(n7702), .C0(
        n4062), .Y(n4061) );
  BUFX4 U11090 ( .A(n7742), .Y(n7752) );
  INVX3 U11091 ( .A(n8275), .Y(n8269) );
  CLKBUFX3 U11092 ( .A(n8173), .Y(n8175) );
  CLKBUFX3 U11093 ( .A(n1749), .Y(n8173) );
  CLKBUFX3 U11094 ( .A(n1751), .Y(n8171) );
  CLKBUFX3 U11095 ( .A(n7732), .Y(n7728) );
  CLKBUFX3 U11096 ( .A(n2655), .Y(n7447) );
  NAND2X1 U11097 ( .A(n4186), .B(n4187), .Y(n2655) );
  AOI222XL U11098 ( .A0(N34766), .A1(n7764), .B0(N32718), .B1(n7704), .C0(
        N31950), .C1(n7761), .Y(n4186) );
  AOI221XL U11099 ( .A0(N33678), .A1(n7872), .B0(N31374), .B1(n7701), .C0(
        n4188), .Y(n4187) );
  CLKBUFX3 U11100 ( .A(n2653), .Y(n7449) );
  NAND2X1 U11101 ( .A(n4168), .B(n4169), .Y(n2653) );
  AOI222XL U11102 ( .A0(N34767), .A1(n7764), .B0(N32719), .B1(n7706), .C0(
        N31951), .C1(n7762), .Y(n4168) );
  AOI221XL U11103 ( .A0(N33679), .A1(n7872), .B0(N31375), .B1(n7702), .C0(
        n4170), .Y(n4169) );
  CLKBUFX3 U11104 ( .A(n2651), .Y(n7451) );
  NAND2X1 U11105 ( .A(n4150), .B(n4151), .Y(n2651) );
  AOI222XL U11106 ( .A0(N34768), .A1(n7764), .B0(N32720), .B1(n7704), .C0(
        N31952), .C1(n7762), .Y(n4150) );
  AOI221XL U11107 ( .A0(N33680), .A1(n7872), .B0(N31376), .B1(n7702), .C0(
        n4152), .Y(n4151) );
  CLKBUFX3 U11108 ( .A(n2649), .Y(n7453) );
  NAND2X1 U11109 ( .A(n4132), .B(n4133), .Y(n2649) );
  AOI222XL U11110 ( .A0(N34769), .A1(n7764), .B0(N32721), .B1(n7706), .C0(
        N31953), .C1(n7762), .Y(n4132) );
  AOI221XL U11111 ( .A0(N33681), .A1(n7872), .B0(N31377), .B1(n7702), .C0(
        n4134), .Y(n4133) );
  CLKBUFX3 U11112 ( .A(n2647), .Y(n7455) );
  NAND2X1 U11113 ( .A(n4114), .B(n4115), .Y(n2647) );
  AOI222XL U11114 ( .A0(N34770), .A1(n3700), .B0(N32722), .B1(n7706), .C0(
        N31954), .C1(n7762), .Y(n4114) );
  AOI221XL U11115 ( .A0(N33682), .A1(n7872), .B0(N31378), .B1(n7702), .C0(
        n4116), .Y(n4115) );
  BUFX4 U11116 ( .A(n7741), .Y(n7751) );
  INVX3 U11117 ( .A(n8329), .Y(n8321) );
  CLKBUFX3 U11118 ( .A(n2663), .Y(n7439) );
  NAND2X1 U11119 ( .A(n4258), .B(n4259), .Y(n2663) );
  AOI222XL U11120 ( .A0(N34762), .A1(n7764), .B0(N32714), .B1(n7705), .C0(
        N31946), .C1(n7763), .Y(n4258) );
  AOI221XL U11121 ( .A0(N33674), .A1(n7872), .B0(N31370), .B1(n7701), .C0(
        n4260), .Y(n4259) );
  CLKBUFX3 U11122 ( .A(n2661), .Y(n7441) );
  NAND2X1 U11123 ( .A(n4240), .B(n4241), .Y(n2661) );
  AOI222XL U11124 ( .A0(N34763), .A1(n7764), .B0(N32715), .B1(n7704), .C0(
        N31947), .C1(n7762), .Y(n4240) );
  AOI221XL U11125 ( .A0(N33675), .A1(n7872), .B0(N31371), .B1(n7701), .C0(
        n4242), .Y(n4241) );
  CLKBUFX3 U11126 ( .A(n2659), .Y(n7443) );
  NAND2X1 U11127 ( .A(n4222), .B(n4223), .Y(n2659) );
  AOI222XL U11128 ( .A0(N34764), .A1(n7764), .B0(N32716), .B1(n7705), .C0(
        N31948), .C1(n7763), .Y(n4222) );
  AOI221XL U11129 ( .A0(N33676), .A1(n7872), .B0(N31372), .B1(n7701), .C0(
        n4224), .Y(n4223) );
  CLKBUFX3 U11130 ( .A(n2657), .Y(n7445) );
  NAND2X1 U11131 ( .A(n4204), .B(n4205), .Y(n2657) );
  AOI222XL U11132 ( .A0(N34765), .A1(n7764), .B0(N32717), .B1(n7704), .C0(
        N31949), .C1(n7762), .Y(n4204) );
  AOI221XL U11133 ( .A0(N33677), .A1(n7872), .B0(N31373), .B1(n7701), .C0(
        n4206), .Y(n4205) );
  INVX3 U11134 ( .A(n8274), .Y(n8271) );
  CLKBUFX3 U11135 ( .A(n7733), .Y(n7726) );
  CLKBUFX3 U11136 ( .A(n7735), .Y(n7722) );
  CLKBUFX3 U11137 ( .A(n7739), .Y(n7714) );
  CLKBUFX3 U11138 ( .A(n7740), .Y(n7712) );
  CLKBUFX3 U11139 ( .A(n2665), .Y(n7437) );
  NAND2X1 U11140 ( .A(n4276), .B(n4277), .Y(n2665) );
  AOI222XL U11141 ( .A0(N34761), .A1(n7764), .B0(N32713), .B1(n8857), .C0(
        N31945), .C1(n7761), .Y(n4276) );
  AOI221XL U11142 ( .A0(N33673), .A1(n7873), .B0(N31369), .B1(n7701), .C0(
        n4278), .Y(n4277) );
  CLKBUFX3 U11143 ( .A(n2671), .Y(n7431) );
  NAND2X1 U11144 ( .A(n4330), .B(n4331), .Y(n2671) );
  AOI222XL U11145 ( .A0(N34758), .A1(n7764), .B0(N32710), .B1(n7705), .C0(
        N31942), .C1(n7762), .Y(n4330) );
  AOI221XL U11146 ( .A0(N33670), .A1(n7873), .B0(N31366), .B1(n7701), .C0(
        n4332), .Y(n4331) );
  CLKBUFX3 U11147 ( .A(n2669), .Y(n7433) );
  NAND2X1 U11148 ( .A(n4312), .B(n4313), .Y(n2669) );
  AOI222XL U11149 ( .A0(N34759), .A1(n7764), .B0(N32711), .B1(n7705), .C0(
        N31943), .C1(n7762), .Y(n4312) );
  AOI221XL U11150 ( .A0(N33671), .A1(n7872), .B0(N31367), .B1(n7701), .C0(
        n4314), .Y(n4313) );
  CLKBUFX3 U11151 ( .A(n2667), .Y(n7435) );
  NAND2X1 U11152 ( .A(n4294), .B(n4295), .Y(n2667) );
  AOI222XL U11153 ( .A0(N34760), .A1(n7764), .B0(N32712), .B1(n7704), .C0(
        N31944), .C1(n7762), .Y(n4294) );
  AOI221XL U11154 ( .A0(N33672), .A1(n7872), .B0(N31368), .B1(n7701), .C0(
        n4296), .Y(n4295) );
  CLKBUFX3 U11155 ( .A(n2679), .Y(n7423) );
  NAND2X1 U11156 ( .A(n4402), .B(n4403), .Y(n2679) );
  AOI222XL U11157 ( .A0(N34754), .A1(n7765), .B0(N32706), .B1(n7705), .C0(
        N31938), .C1(n7763), .Y(n4402) );
  AOI221XL U11158 ( .A0(N33666), .A1(n7873), .B0(N31362), .B1(n7701), .C0(
        n4404), .Y(n4403) );
  CLKBUFX3 U11159 ( .A(n2677), .Y(n7425) );
  NAND2X1 U11160 ( .A(n4384), .B(n4385), .Y(n2677) );
  AOI222XL U11161 ( .A0(N34755), .A1(n7765), .B0(N32707), .B1(n7705), .C0(
        N31939), .C1(n7762), .Y(n4384) );
  AOI221XL U11162 ( .A0(N33667), .A1(n7873), .B0(N31363), .B1(n7701), .C0(
        n4386), .Y(n4385) );
  CLKBUFX3 U11163 ( .A(n2675), .Y(n7427) );
  NAND2X1 U11164 ( .A(n4366), .B(n4367), .Y(n2675) );
  AOI222XL U11165 ( .A0(N34756), .A1(n7765), .B0(N32708), .B1(n7705), .C0(
        N31940), .C1(n7762), .Y(n4366) );
  AOI221XL U11166 ( .A0(N33668), .A1(n7872), .B0(N31364), .B1(n7701), .C0(
        n4368), .Y(n4367) );
  CLKBUFX3 U11167 ( .A(n2673), .Y(n7429) );
  NAND2X1 U11168 ( .A(n4348), .B(n4349), .Y(n2673) );
  AOI222XL U11169 ( .A0(N34757), .A1(n7765), .B0(N32709), .B1(n7705), .C0(
        N31941), .C1(n7762), .Y(n4348) );
  AOI221XL U11170 ( .A0(N33669), .A1(n7872), .B0(N31365), .B1(n7701), .C0(
        n4350), .Y(n4349) );
  CLKBUFX3 U11171 ( .A(n7737), .Y(n7717) );
  CLKBUFX3 U11172 ( .A(n2683), .Y(n7419) );
  NAND2X1 U11173 ( .A(n4438), .B(n4439), .Y(n2683) );
  AOI222XL U11174 ( .A0(N34752), .A1(n7765), .B0(N32704), .B1(n7705), .C0(
        N31936), .C1(n8860), .Y(n4438) );
  AOI221XL U11175 ( .A0(N33664), .A1(n7873), .B0(N31360), .B1(n7701), .C0(
        n4440), .Y(n4439) );
  CLKBUFX3 U11176 ( .A(n2685), .Y(n7417) );
  NAND2X1 U11177 ( .A(n4456), .B(n4457), .Y(n2685) );
  AOI222XL U11178 ( .A0(N34751), .A1(n7765), .B0(N32703), .B1(n7705), .C0(
        N31935), .C1(n7761), .Y(n4456) );
  AOI221XL U11179 ( .A0(N33663), .A1(n7873), .B0(N31359), .B1(n7701), .C0(
        n4458), .Y(n4457) );
  CLKBUFX3 U11180 ( .A(n2681), .Y(n7421) );
  NAND2X1 U11181 ( .A(n4420), .B(n4421), .Y(n2681) );
  AOI222XL U11182 ( .A0(N34753), .A1(n7765), .B0(N32705), .B1(n7705), .C0(
        N31937), .C1(n7763), .Y(n4420) );
  AOI221XL U11183 ( .A0(N33665), .A1(n7873), .B0(N31361), .B1(n7701), .C0(
        n4422), .Y(n4421) );
  CLKBUFX3 U11184 ( .A(n2697), .Y(n7405) );
  NAND2X1 U11185 ( .A(n4564), .B(n4565), .Y(n2697) );
  AOI222XL U11186 ( .A0(N34745), .A1(n7766), .B0(N32697), .B1(n7705), .C0(
        N31929), .C1(n8860), .Y(n4564) );
  AOI221XL U11187 ( .A0(N33657), .A1(n7873), .B0(N31353), .B1(n7700), .C0(
        n4566), .Y(n4565) );
  CLKBUFX3 U11188 ( .A(n2695), .Y(n7407) );
  NAND2X1 U11189 ( .A(n4546), .B(n4547), .Y(n2695) );
  AOI222XL U11190 ( .A0(N34746), .A1(n7765), .B0(N32698), .B1(n7705), .C0(
        N31930), .C1(n7763), .Y(n4546) );
  AOI221XL U11191 ( .A0(N33658), .A1(n7874), .B0(N31354), .B1(n7700), .C0(
        n4548), .Y(n4547) );
  CLKBUFX3 U11192 ( .A(n2693), .Y(n7409) );
  NAND2X1 U11193 ( .A(n4528), .B(n4529), .Y(n2693) );
  AOI222XL U11194 ( .A0(N34747), .A1(n7765), .B0(N32699), .B1(n7705), .C0(
        N31931), .C1(n7761), .Y(n4528) );
  AOI221XL U11195 ( .A0(N33659), .A1(n7874), .B0(N31355), .B1(n7701), .C0(
        n4530), .Y(n4529) );
  CLKBUFX3 U11196 ( .A(n2691), .Y(n7411) );
  NAND2X1 U11197 ( .A(n4510), .B(n4511), .Y(n2691) );
  AOI222XL U11198 ( .A0(N34748), .A1(n7765), .B0(N32700), .B1(n7705), .C0(
        N31932), .C1(n7763), .Y(n4510) );
  AOI221XL U11199 ( .A0(N33660), .A1(n7873), .B0(N31356), .B1(n7701), .C0(
        n4512), .Y(n4511) );
  CLKBUFX3 U11200 ( .A(n2689), .Y(n7413) );
  NAND2X1 U11201 ( .A(n4492), .B(n4493), .Y(n2689) );
  AOI222XL U11202 ( .A0(N34749), .A1(n7765), .B0(N32701), .B1(n7705), .C0(
        N31933), .C1(n7761), .Y(n4492) );
  AOI221XL U11203 ( .A0(N33661), .A1(n7873), .B0(N31357), .B1(n7701), .C0(
        n4494), .Y(n4493) );
  CLKBUFX3 U11204 ( .A(n2687), .Y(n7415) );
  NAND2X1 U11205 ( .A(n4474), .B(n4475), .Y(n2687) );
  AOI222XL U11206 ( .A0(N34750), .A1(n7765), .B0(N32702), .B1(n7705), .C0(
        N31934), .C1(n7761), .Y(n4474) );
  AOI221XL U11207 ( .A0(N33662), .A1(n7873), .B0(N31358), .B1(n7701), .C0(
        n4476), .Y(n4475) );
  CLKBUFX3 U11208 ( .A(n7731), .Y(n7730) );
  CLKBUFX3 U11209 ( .A(n1751), .Y(n8170) );
  CLKBUFX3 U11210 ( .A(n2703), .Y(n7399) );
  NAND2X1 U11211 ( .A(n4618), .B(n4619), .Y(n2703) );
  AOI222XL U11212 ( .A0(N34742), .A1(n7766), .B0(N32694), .B1(n7704), .C0(
        N31926), .C1(n8860), .Y(n4618) );
  AOI221XL U11213 ( .A0(N33654), .A1(n7874), .B0(N31350), .B1(n7700), .C0(
        n4620), .Y(n4619) );
  CLKBUFX3 U11214 ( .A(n2701), .Y(n7401) );
  NAND2X1 U11215 ( .A(n4600), .B(n4601), .Y(n2701) );
  AOI222XL U11216 ( .A0(N34743), .A1(n7766), .B0(N32695), .B1(n7704), .C0(
        N31927), .C1(n7761), .Y(n4600) );
  AOI221XL U11217 ( .A0(N33655), .A1(n7874), .B0(N31351), .B1(n7701), .C0(
        n4602), .Y(n4601) );
  CLKBUFX3 U11218 ( .A(n2699), .Y(n7403) );
  NAND2X1 U11219 ( .A(n4582), .B(n4583), .Y(n2699) );
  AOI222XL U11220 ( .A0(N34744), .A1(n7766), .B0(N32696), .B1(n7705), .C0(
        N31928), .C1(n8860), .Y(n4582) );
  AOI221XL U11221 ( .A0(N33656), .A1(n7873), .B0(N31352), .B1(n7700), .C0(
        n4584), .Y(n4583) );
  CLKBUFX3 U11222 ( .A(n8771), .Y(n7505) );
  CLKINVX1 U11223 ( .A(N25659), .Y(n8771) );
  CLKBUFX3 U11224 ( .A(n8770), .Y(n7504) );
  CLKINVX1 U11225 ( .A(N25660), .Y(n8770) );
  CLKBUFX3 U11226 ( .A(n8768), .Y(n7564) );
  CLKBUFX3 U11227 ( .A(n8768), .Y(n7565) );
  CLKBUFX3 U11228 ( .A(n8768), .Y(n7566) );
  CLKBUFX3 U11229 ( .A(n2705), .Y(n7397) );
  NAND2X1 U11230 ( .A(n4636), .B(n4637), .Y(n2705) );
  AOI222XL U11231 ( .A0(N34741), .A1(n7766), .B0(N32693), .B1(n7704), .C0(
        N31925), .C1(n7761), .Y(n4636) );
  AOI221XL U11232 ( .A0(N33653), .A1(n7874), .B0(N31349), .B1(n7700), .C0(
        n4638), .Y(n4637) );
  CLKBUFX3 U11233 ( .A(n2711), .Y(n7391) );
  NAND2X1 U11234 ( .A(n4690), .B(n4691), .Y(n2711) );
  AOI222XL U11235 ( .A0(N34738), .A1(n7766), .B0(N32690), .B1(n7704), .C0(
        N31922), .C1(n7761), .Y(n4690) );
  AOI221XL U11236 ( .A0(N33650), .A1(n7874), .B0(N31346), .B1(n7700), .C0(
        n4692), .Y(n4691) );
  CLKBUFX3 U11237 ( .A(n2709), .Y(n7393) );
  NAND2X1 U11238 ( .A(n4672), .B(n4673), .Y(n2709) );
  AOI222XL U11239 ( .A0(N34739), .A1(n7766), .B0(N32691), .B1(n7704), .C0(
        N31923), .C1(n7761), .Y(n4672) );
  AOI221XL U11240 ( .A0(N33651), .A1(n7874), .B0(N31347), .B1(n7700), .C0(
        n4674), .Y(n4673) );
  CLKBUFX3 U11241 ( .A(n2707), .Y(n7395) );
  NAND2X1 U11242 ( .A(n4654), .B(n4655), .Y(n2707) );
  AOI222XL U11243 ( .A0(N34740), .A1(n7766), .B0(N32692), .B1(n7704), .C0(
        N31924), .C1(n7761), .Y(n4654) );
  AOI221XL U11244 ( .A0(N33652), .A1(n7874), .B0(N31348), .B1(n7700), .C0(
        n4656), .Y(n4655) );
  CLKBUFX3 U11245 ( .A(n8774), .Y(n7508) );
  CLKINVX1 U11246 ( .A(N25656), .Y(n8774) );
  CLKBUFX3 U11247 ( .A(n8773), .Y(n7507) );
  CLKINVX1 U11248 ( .A(N25657), .Y(n8773) );
  CLKBUFX3 U11249 ( .A(n8772), .Y(n7506) );
  CLKINVX1 U11250 ( .A(N25658), .Y(n8772) );
  CLKBUFX3 U11251 ( .A(n7731), .Y(n7729) );
  CLKBUFX3 U11252 ( .A(n7733), .Y(n7725) );
  CLKBUFX3 U11253 ( .A(n7740), .Y(n7713) );
  CLKBUFX3 U11254 ( .A(n2723), .Y(n7379) );
  NAND2X1 U11255 ( .A(n4798), .B(n4799), .Y(n2723) );
  AOI222XL U11256 ( .A0(N34732), .A1(n7764), .B0(N32684), .B1(n7704), .C0(
        N31916), .C1(n7761), .Y(n4798) );
  AOI221XL U11257 ( .A0(N33644), .A1(n7875), .B0(N31340), .B1(n7700), .C0(
        n4800), .Y(n4799) );
  CLKBUFX3 U11258 ( .A(n2721), .Y(n7381) );
  NAND2X1 U11259 ( .A(n4780), .B(n4781), .Y(n2721) );
  AOI222XL U11260 ( .A0(N34733), .A1(n7764), .B0(N32685), .B1(n7704), .C0(
        N31917), .C1(n7761), .Y(n4780) );
  AOI221XL U11261 ( .A0(N33645), .A1(n7874), .B0(N31341), .B1(n7700), .C0(
        n4782), .Y(n4781) );
  CLKBUFX3 U11262 ( .A(n2719), .Y(n7383) );
  NAND2X1 U11263 ( .A(n4762), .B(n4763), .Y(n2719) );
  AOI222XL U11264 ( .A0(N34734), .A1(n7766), .B0(N32686), .B1(n7704), .C0(
        N31918), .C1(n7761), .Y(n4762) );
  AOI221XL U11265 ( .A0(N33646), .A1(n7874), .B0(N31342), .B1(n7700), .C0(
        n4764), .Y(n4763) );
  CLKBUFX3 U11266 ( .A(n2717), .Y(n7385) );
  NAND2X1 U11267 ( .A(n4744), .B(n4745), .Y(n2717) );
  AOI222XL U11268 ( .A0(N34735), .A1(n7766), .B0(N32687), .B1(n7704), .C0(
        N31919), .C1(n7761), .Y(n4744) );
  AOI221XL U11269 ( .A0(N33647), .A1(n7874), .B0(N31343), .B1(n7700), .C0(
        n4746), .Y(n4745) );
  CLKBUFX3 U11270 ( .A(n2715), .Y(n7387) );
  NAND2X1 U11271 ( .A(n4726), .B(n4727), .Y(n2715) );
  AOI222XL U11272 ( .A0(N34736), .A1(n7766), .B0(N32688), .B1(n7704), .C0(
        N31920), .C1(n7761), .Y(n4726) );
  AOI221XL U11273 ( .A0(N33648), .A1(n7874), .B0(N31344), .B1(n7700), .C0(
        n4728), .Y(n4727) );
  CLKBUFX3 U11274 ( .A(n2713), .Y(n7389) );
  NAND2X1 U11275 ( .A(n4708), .B(n4709), .Y(n2713) );
  AOI222XL U11276 ( .A0(N34737), .A1(n7766), .B0(N32689), .B1(n7704), .C0(
        N31921), .C1(n7761), .Y(n4708) );
  AOI221XL U11277 ( .A0(N33649), .A1(n7874), .B0(N31345), .B1(n7700), .C0(
        n4710), .Y(n4709) );
  CLKBUFX3 U11278 ( .A(n8777), .Y(n7511) );
  CLKINVX1 U11279 ( .A(N25653), .Y(n8777) );
  CLKBUFX3 U11280 ( .A(n8776), .Y(n7510) );
  CLKINVX1 U11281 ( .A(N25654), .Y(n8776) );
  CLKBUFX3 U11282 ( .A(n8775), .Y(n7509) );
  CLKINVX1 U11283 ( .A(N25655), .Y(n8775) );
  CLKBUFX3 U11284 ( .A(n7712), .Y(n7721) );
  CLKBUFX3 U11285 ( .A(n2725), .Y(n7377) );
  NAND2X1 U11286 ( .A(n4816), .B(n4817), .Y(n2725) );
  AOI222XL U11287 ( .A0(N34731), .A1(n7765), .B0(N32683), .B1(n7704), .C0(
        N31915), .C1(n7761), .Y(n4816) );
  AOI221XL U11288 ( .A0(N33643), .A1(n7875), .B0(N31339), .B1(n7700), .C0(
        n4818), .Y(n4817) );
  CLKBUFX3 U11289 ( .A(n2727), .Y(n7375) );
  NAND2X1 U11290 ( .A(n4870), .B(n4871), .Y(n2727) );
  AOI222XL U11291 ( .A0(N34730), .A1(n7765), .B0(N32682), .B1(n7704), .C0(
        N31914), .C1(n7763), .Y(n4870) );
  AOI221XL U11292 ( .A0(N33642), .A1(n7875), .B0(N31338), .B1(n7700), .C0(
        n4872), .Y(n4871) );
  CLKBUFX3 U11293 ( .A(n8780), .Y(n7514) );
  CLKINVX1 U11294 ( .A(N25650), .Y(n8780) );
  CLKBUFX3 U11295 ( .A(n8779), .Y(n7513) );
  CLKINVX1 U11296 ( .A(N25651), .Y(n8779) );
  CLKBUFX3 U11297 ( .A(n8778), .Y(n7512) );
  CLKINVX1 U11298 ( .A(N25652), .Y(n8778) );
  CLKBUFX3 U11299 ( .A(n8783), .Y(n7517) );
  CLKINVX1 U11300 ( .A(N25647), .Y(n8783) );
  CLKBUFX3 U11301 ( .A(n8782), .Y(n7516) );
  CLKINVX1 U11302 ( .A(N25648), .Y(n8782) );
  CLKBUFX3 U11303 ( .A(n8781), .Y(n7515) );
  CLKINVX1 U11304 ( .A(N25649), .Y(n8781) );
  CLKBUFX3 U11305 ( .A(n6979), .Y(n6986) );
  CLKBUFX3 U11306 ( .A(n8786), .Y(n7520) );
  CLKINVX1 U11307 ( .A(N25644), .Y(n8786) );
  CLKBUFX3 U11308 ( .A(n8785), .Y(n7519) );
  CLKINVX1 U11309 ( .A(N25645), .Y(n8785) );
  CLKBUFX3 U11310 ( .A(n8784), .Y(n7518) );
  CLKINVX1 U11311 ( .A(N25646), .Y(n8784) );
  CLKBUFX3 U11312 ( .A(n7202), .Y(n7209) );
  CLKBUFX3 U11313 ( .A(n6979), .Y(n6987) );
  CLKBUFX3 U11314 ( .A(n8788), .Y(n7522) );
  CLKINVX1 U11315 ( .A(N25642), .Y(n8788) );
  CLKBUFX3 U11316 ( .A(n8787), .Y(n7521) );
  CLKINVX1 U11317 ( .A(N25643), .Y(n8787) );
  CLKBUFX3 U11318 ( .A(n7214), .Y(n7221) );
  CLKBUFX3 U11319 ( .A(n6994), .Y(n7000) );
  CLKBUFX3 U11320 ( .A(n8791), .Y(n7525) );
  CLKINVX1 U11321 ( .A(N25639), .Y(n8791) );
  CLKBUFX3 U11322 ( .A(n8790), .Y(n7524) );
  CLKINVX1 U11323 ( .A(N25640), .Y(n8790) );
  CLKBUFX3 U11324 ( .A(n8789), .Y(n7523) );
  CLKINVX1 U11325 ( .A(N25641), .Y(n8789) );
  CLKBUFX3 U11326 ( .A(n6978), .Y(n6988) );
  CLKBUFX3 U11327 ( .A(n8794), .Y(n7528) );
  CLKINVX1 U11328 ( .A(N25636), .Y(n8794) );
  CLKBUFX3 U11329 ( .A(n8793), .Y(n7527) );
  CLKINVX1 U11330 ( .A(N25637), .Y(n8793) );
  CLKBUFX3 U11331 ( .A(n8792), .Y(n7526) );
  CLKINVX1 U11332 ( .A(N25638), .Y(n8792) );
  CLKBUFX3 U11333 ( .A(n8797), .Y(n7531) );
  CLKINVX1 U11334 ( .A(N25633), .Y(n8797) );
  CLKBUFX3 U11335 ( .A(n8796), .Y(n7530) );
  CLKINVX1 U11336 ( .A(N25634), .Y(n8796) );
  CLKBUFX3 U11337 ( .A(n8795), .Y(n7529) );
  CLKINVX1 U11338 ( .A(N25635), .Y(n8795) );
  CLKBUFX3 U11339 ( .A(n7740), .Y(n7720) );
  CLKBUFX3 U11340 ( .A(n8800), .Y(n7534) );
  CLKINVX1 U11341 ( .A(N25630), .Y(n8800) );
  CLKBUFX3 U11342 ( .A(n8799), .Y(n7533) );
  CLKINVX1 U11343 ( .A(N25631), .Y(n8799) );
  CLKBUFX3 U11344 ( .A(n8798), .Y(n7532) );
  CLKINVX1 U11345 ( .A(N25632), .Y(n8798) );
  CLKBUFX3 U11346 ( .A(n8803), .Y(n7537) );
  CLKINVX1 U11347 ( .A(N25627), .Y(n8803) );
  CLKBUFX3 U11348 ( .A(n8802), .Y(n7536) );
  CLKINVX1 U11349 ( .A(N25628), .Y(n8802) );
  CLKBUFX3 U11350 ( .A(n8801), .Y(n7535) );
  CLKINVX1 U11351 ( .A(N25629), .Y(n8801) );
  CLKBUFX3 U11352 ( .A(n8805), .Y(n7539) );
  CLKINVX1 U11353 ( .A(N25625), .Y(n8805) );
  CLKBUFX3 U11354 ( .A(n8804), .Y(n7538) );
  CLKINVX1 U11355 ( .A(N25626), .Y(n8804) );
  CLKBUFX3 U11356 ( .A(n8808), .Y(n7542) );
  CLKINVX1 U11357 ( .A(N25622), .Y(n8808) );
  CLKBUFX3 U11358 ( .A(n8807), .Y(n7541) );
  CLKINVX1 U11359 ( .A(N25623), .Y(n8807) );
  CLKBUFX3 U11360 ( .A(n8806), .Y(n7540) );
  CLKINVX1 U11361 ( .A(N25624), .Y(n8806) );
  CLKBUFX3 U11362 ( .A(n8811), .Y(n7545) );
  CLKINVX1 U11363 ( .A(N25619), .Y(n8811) );
  CLKBUFX3 U11364 ( .A(n8810), .Y(n7544) );
  CLKINVX1 U11365 ( .A(N25620), .Y(n8810) );
  CLKBUFX3 U11366 ( .A(n8809), .Y(n7543) );
  CLKINVX1 U11367 ( .A(N25621), .Y(n8809) );
  CLKBUFX3 U11368 ( .A(n8814), .Y(n7548) );
  CLKINVX1 U11369 ( .A(N25616), .Y(n8814) );
  CLKBUFX3 U11370 ( .A(n8813), .Y(n7547) );
  CLKINVX1 U11371 ( .A(N25617), .Y(n8813) );
  CLKBUFX3 U11372 ( .A(n8812), .Y(n7546) );
  CLKINVX1 U11373 ( .A(N25618), .Y(n8812) );
  CLKBUFX3 U11374 ( .A(n8817), .Y(n7551) );
  CLKINVX1 U11375 ( .A(N25613), .Y(n8817) );
  CLKBUFX3 U11376 ( .A(n8816), .Y(n7550) );
  CLKINVX1 U11377 ( .A(N25614), .Y(n8816) );
  CLKBUFX3 U11378 ( .A(n8815), .Y(n7549) );
  CLKINVX1 U11379 ( .A(N25615), .Y(n8815) );
  CLKBUFX3 U11380 ( .A(n8820), .Y(n7554) );
  CLKINVX1 U11381 ( .A(N25610), .Y(n8820) );
  CLKBUFX3 U11382 ( .A(n8819), .Y(n7553) );
  CLKINVX1 U11383 ( .A(N25611), .Y(n8819) );
  CLKBUFX3 U11384 ( .A(n8818), .Y(n7552) );
  CLKINVX1 U11385 ( .A(N25612), .Y(n8818) );
  CLKBUFX3 U11386 ( .A(n8822), .Y(n7556) );
  CLKINVX1 U11387 ( .A(N25608), .Y(n8822) );
  CLKBUFX3 U11388 ( .A(n8821), .Y(n7555) );
  CLKINVX1 U11389 ( .A(N25609), .Y(n8821) );
  CLKBUFX3 U11390 ( .A(n8825), .Y(n7559) );
  CLKINVX1 U11391 ( .A(N25605), .Y(n8825) );
  CLKBUFX3 U11392 ( .A(n8824), .Y(n7558) );
  CLKINVX1 U11393 ( .A(N25606), .Y(n8824) );
  CLKBUFX3 U11394 ( .A(n8823), .Y(n7557) );
  CLKINVX1 U11395 ( .A(N25607), .Y(n8823) );
  CLKBUFX3 U11396 ( .A(n8828), .Y(n7562) );
  CLKINVX1 U11397 ( .A(N25602), .Y(n8828) );
  CLKBUFX3 U11398 ( .A(n8827), .Y(n7561) );
  CLKINVX1 U11399 ( .A(N25603), .Y(n8827) );
  CLKBUFX3 U11400 ( .A(n8826), .Y(n7560) );
  CLKINVX1 U11401 ( .A(N25604), .Y(n8826) );
  CLKBUFX3 U11402 ( .A(n8829), .Y(n7563) );
  CLKINVX1 U11403 ( .A(N25601), .Y(n8829) );
  CLKBUFX3 U11404 ( .A(n8122), .Y(n8125) );
  CLKBUFX3 U11405 ( .A(n8045), .Y(n8048) );
  CLKBUFX3 U11406 ( .A(n8122), .Y(n8124) );
  CLKBUFX3 U11407 ( .A(n3652), .Y(n7970) );
  CLKBUFX3 U11408 ( .A(n8045), .Y(n8047) );
  CLKBUFX3 U11409 ( .A(n8096), .Y(n8099) );
  CLKBUFX3 U11410 ( .A(n3652), .Y(n7969) );
  CLKBUFX3 U11411 ( .A(n8096), .Y(n8098) );
  CLKBUFX3 U11412 ( .A(n8122), .Y(n8123) );
  CLKBUFX3 U11413 ( .A(n2601), .Y(n8134) );
  CLKBUFX3 U11414 ( .A(n3154), .Y(n8057) );
  CLKBUFX3 U11415 ( .A(n3154), .Y(n8056) );
  CLKBUFX3 U11416 ( .A(n2601), .Y(n8133) );
  CLKBUFX3 U11417 ( .A(n3154), .Y(n8055) );
  CLKBUFX3 U11418 ( .A(n2601), .Y(n8132) );
  CLKBUFX3 U11419 ( .A(n3362), .Y(n8026) );
  CLKBUFX3 U11420 ( .A(n3010), .Y(n8090) );
  CLKBUFX3 U11421 ( .A(n7988), .Y(n7989) );
  CLKBUFX3 U11422 ( .A(n8052), .Y(n8053) );
  CLKBUFX3 U11423 ( .A(n8103), .Y(n8104) );
  CLKBUFX3 U11424 ( .A(n8116), .Y(n8117) );
  CLKBUFX3 U11425 ( .A(n6609), .Y(n8129) );
  CLKBUFX3 U11426 ( .A(n3226), .Y(n8044) );
  CLKBUFX3 U11427 ( .A(n2943), .Y(n8095) );
  CLKBUFX3 U11428 ( .A(n2736), .Y(n8121) );
  CLKBUFX3 U11429 ( .A(n3654), .Y(n7968) );
  CLKBUFX3 U11430 ( .A(n3226), .Y(n8043) );
  CLKBUFX3 U11431 ( .A(n2943), .Y(n8094) );
  CLKBUFX3 U11432 ( .A(n2736), .Y(n8120) );
  CLKBUFX3 U11433 ( .A(n3654), .Y(n7967) );
  CLKBUFX3 U11434 ( .A(n3226), .Y(n8042) );
  CLKBUFX3 U11435 ( .A(n2943), .Y(n8093) );
  CLKBUFX3 U11436 ( .A(n2736), .Y(n8119) );
  CLKBUFX3 U11437 ( .A(n3654), .Y(n7966) );
  AND2X2 U11438 ( .A(n7973), .B(n3649), .Y(n4821) );
  CLKBUFX3 U11439 ( .A(n8110), .Y(n8109) );
  CLKBUFX3 U11440 ( .A(n3431), .Y(n8013) );
  CLKBUFX3 U11441 ( .A(n3362), .Y(n8027) );
  CLKBUFX3 U11442 ( .A(n8039), .Y(n8040) );
  CLKBUFX3 U11443 ( .A(n3081), .Y(n8077) );
  CLKBUFX3 U11444 ( .A(n3010), .Y(n8091) );
  CLKBUFX3 U11445 ( .A(n8013), .Y(n8014) );
  CLKBUFX3 U11446 ( .A(n8077), .Y(n8078) );
  CLKBUFX3 U11447 ( .A(n8169), .Y(n8167) );
  CLKBUFX3 U11448 ( .A(n8003), .Y(n8002) );
  CLKBUFX3 U11449 ( .A(n8013), .Y(n8015) );
  CLKBUFX3 U11450 ( .A(n8077), .Y(n8079) );
  CLKBUFX3 U11451 ( .A(n8091), .Y(n8092) );
  CLKBUFX3 U11452 ( .A(n8156), .Y(n8155) );
  CLKBUFX3 U11453 ( .A(n8169), .Y(n8168) );
  CLKBUFX3 U11454 ( .A(n8064), .Y(n8065) );
  CLKBUFX3 U11455 ( .A(n6609), .Y(n8130) );
  CLKBUFX3 U11456 ( .A(n8141), .Y(n8142) );
  CLKBUFX3 U11457 ( .A(n8052), .Y(n8054) );
  CLKBUFX3 U11458 ( .A(n8065), .Y(n8066) );
  CLKBUFX3 U11459 ( .A(n8117), .Y(n8118) );
  CLKBUFX3 U11460 ( .A(n8142), .Y(n8143) );
  CLKBUFX3 U11461 ( .A(n7989), .Y(n7990) );
  CLKBUFX3 U11462 ( .A(n7886), .Y(n7881) );
  CLKBUFX3 U11463 ( .A(n7991), .Y(n7992) );
  CLKBUFX3 U11464 ( .A(n2595), .Y(n8144) );
  CLKINVX1 U11465 ( .A(n4853), .Y(n8848) );
  CLKBUFX3 U11466 ( .A(n3662), .Y(n7958) );
  CLKBUFX3 U11467 ( .A(n3662), .Y(n7957) );
  CLKBUFX3 U11468 ( .A(n3662), .Y(n7956) );
  CLKBUFX3 U11469 ( .A(n3498), .Y(n8006) );
  CLKBUFX3 U11470 ( .A(n3676), .Y(n7931) );
  CLKBUFX3 U11471 ( .A(n7929), .Y(n7930) );
  CLKBUFX3 U11472 ( .A(n3700), .Y(n7766) );
  CLKBUFX3 U11473 ( .A(n3700), .Y(n7765) );
  CLKBUFX3 U11474 ( .A(n3700), .Y(n7764) );
  CLKBUFX3 U11475 ( .A(n3665), .Y(n7952) );
  CLKBUFX3 U11476 ( .A(n3665), .Y(n7951) );
  CLKBUFX3 U11477 ( .A(n3665), .Y(n7950) );
  CLKBUFX3 U11478 ( .A(n3669), .Y(n7943) );
  CLKBUFX3 U11479 ( .A(n3675), .Y(n7934) );
  CLKBUFX3 U11480 ( .A(n3669), .Y(n7942) );
  CLKBUFX3 U11481 ( .A(n3675), .Y(n7933) );
  CLKBUFX3 U11482 ( .A(n3675), .Y(n7932) );
  CLKBUFX3 U11483 ( .A(n3669), .Y(n7941) );
  CLKBUFX3 U11484 ( .A(n3671), .Y(n7935) );
  CLKBUFX3 U11485 ( .A(n7767), .Y(n7780) );
  CLKBUFX3 U11486 ( .A(n8857), .Y(n7704) );
  CLKBUFX3 U11487 ( .A(n2595), .Y(n8145) );
  CLKBUFX3 U11488 ( .A(n8029), .Y(n8030) );
  CLKBUFX3 U11489 ( .A(n8145), .Y(n8146) );
  CLKBUFX3 U11490 ( .A(n8029), .Y(n8031) );
  CLKBUFX3 U11491 ( .A(n8145), .Y(n8147) );
  CLKBUFX3 U11492 ( .A(n8029), .Y(n8032) );
  CLKBUFX3 U11493 ( .A(n7805), .Y(n7797) );
  CLKBUFX3 U11494 ( .A(n7887), .Y(n7879) );
  CLKBUFX3 U11495 ( .A(n7887), .Y(n7878) );
  CLKBUFX3 U11496 ( .A(n7806), .Y(n7796) );
  CLKBUFX3 U11497 ( .A(n7806), .Y(n7795) );
  CLKBUFX3 U11498 ( .A(n7806), .Y(n7794) );
  CLKBUFX3 U11499 ( .A(n7888), .Y(n7877) );
  CLKBUFX3 U11500 ( .A(n7888), .Y(n7876) );
  CLKBUFX3 U11501 ( .A(n8157), .Y(n8158) );
  CLKBUFX3 U11502 ( .A(n7991), .Y(n7993) );
  CLKBUFX3 U11503 ( .A(n8158), .Y(n8160) );
  CLKBUFX3 U11504 ( .A(n7993), .Y(n7994) );
  CLKBUFX3 U11505 ( .A(n8157), .Y(n8159) );
  CLKBUFX3 U11506 ( .A(n8067), .Y(n8068) );
  CLKBUFX3 U11507 ( .A(n8067), .Y(n8069) );
  CLKBUFX3 U11508 ( .A(n8083), .Y(n8081) );
  CLKBUFX3 U11509 ( .A(n8080), .Y(n8082) );
  CLKBUFX3 U11510 ( .A(n6602), .Y(n8016) );
  CLKBUFX3 U11511 ( .A(n8019), .Y(n8017) );
  CLKBUFX3 U11512 ( .A(n6602), .Y(n8018) );
  CLKBUFX3 U11513 ( .A(n7804), .Y(n7803) );
  CLKBUFX3 U11514 ( .A(n6603), .Y(n7949) );
  CLKBUFX3 U11515 ( .A(n6603), .Y(n7948) );
  CLKBUFX3 U11516 ( .A(n6603), .Y(n7947) );
  CLKBUFX3 U11517 ( .A(n7767), .Y(n7781) );
  CLKBUFX3 U11518 ( .A(n8856), .Y(n7703) );
  CLKBUFX3 U11519 ( .A(n7767), .Y(n7782) );
  CLKBUFX3 U11520 ( .A(n6719), .Y(n7699) );
  CLKBUFX3 U11521 ( .A(n7686), .Y(n7687) );
  CLKBUFX3 U11522 ( .A(n6721), .Y(n7689) );
  CLKBUFX3 U11523 ( .A(n7690), .Y(n7691) );
  CLKBUFX3 U11524 ( .A(n6723), .Y(n7693) );
  CLKBUFX3 U11525 ( .A(n6724), .Y(n7695) );
  CLKBUFX3 U11526 ( .A(n6725), .Y(n7671) );
  CLKBUFX3 U11527 ( .A(n6726), .Y(n7673) );
  CLKBUFX3 U11528 ( .A(n7674), .Y(n7675) );
  CLKBUFX3 U11529 ( .A(n6728), .Y(n7677) );
  CLKBUFX3 U11530 ( .A(n7678), .Y(n7679) );
  CLKBUFX3 U11531 ( .A(n6730), .Y(n7681) );
  CLKBUFX3 U11532 ( .A(n6731), .Y(n7683) );
  CLKBUFX3 U11533 ( .A(n6732), .Y(n7685) );
  CLKBUFX3 U11534 ( .A(n6733), .Y(n7697) );
  CLKBUFX3 U11535 ( .A(n6734), .Y(n7669) );
  CLKBUFX3 U11536 ( .A(n8161), .Y(n8162) );
  CLKBUFX3 U11537 ( .A(n7807), .Y(n7813) );
  CLKBUFX3 U11538 ( .A(n7886), .Y(n7880) );
  INVX3 U11539 ( .A(n7833), .Y(n7831) );
  INVX3 U11540 ( .A(n7852), .Y(n7850) );
  INVX3 U11541 ( .A(n7834), .Y(n7830) );
  INVX3 U11542 ( .A(n7853), .Y(n7849) );
  CLKBUFX3 U11543 ( .A(n8406), .Y(n7361) );
  CLKBUFX3 U11544 ( .A(n8406), .Y(n7362) );
  CLKBUFX3 U11545 ( .A(n8406), .Y(n7363) );
  CLKBUFX3 U11546 ( .A(n8406), .Y(n7364) );
  CLKBUFX3 U11547 ( .A(n8406), .Y(n7365) );
  CLKBUFX3 U11548 ( .A(n8406), .Y(n7366) );
  CLKBUFX3 U11549 ( .A(n7804), .Y(n7802) );
  CLKBUFX3 U11550 ( .A(n7880), .Y(n7885) );
  CLKBUFX3 U11551 ( .A(n7846), .Y(n7835) );
  CLKBUFX3 U11552 ( .A(n7866), .Y(n7854) );
  CLKBUFX3 U11553 ( .A(n7880), .Y(n7884) );
  CLKBUFX3 U11554 ( .A(n7846), .Y(n7836) );
  CLKBUFX3 U11555 ( .A(n7866), .Y(n7855) );
  CLKBUFX3 U11556 ( .A(n7804), .Y(n7801) );
  CLKBUFX3 U11557 ( .A(n7846), .Y(n7837) );
  CLKBUFX3 U11558 ( .A(n7866), .Y(n7856) );
  CLKBUFX3 U11559 ( .A(n7846), .Y(n7838) );
  CLKBUFX3 U11560 ( .A(n7847), .Y(n7857) );
  CLKBUFX3 U11561 ( .A(n7859), .Y(n7858) );
  CLKBUFX3 U11562 ( .A(n7802), .Y(n7800) );
  CLKBUFX3 U11563 ( .A(n7845), .Y(n7839) );
  CLKBUFX3 U11564 ( .A(n7847), .Y(n7859) );
  CLKBUFX3 U11565 ( .A(n7845), .Y(n7840) );
  CLKBUFX3 U11566 ( .A(n7798), .Y(n7799) );
  CLKBUFX3 U11567 ( .A(n7845), .Y(n7841) );
  CLKBUFX3 U11568 ( .A(n7865), .Y(n7860) );
  CLKBUFX3 U11569 ( .A(n7844), .Y(n7842) );
  CLKBUFX3 U11570 ( .A(n7865), .Y(n7861) );
  CLKBUFX3 U11571 ( .A(n7880), .Y(n7883) );
  CLKBUFX3 U11572 ( .A(n7860), .Y(n7862) );
  CLKBUFX3 U11573 ( .A(n7801), .Y(n7798) );
  CLKBUFX3 U11574 ( .A(n7886), .Y(n7882) );
  CLKBUFX3 U11575 ( .A(n7844), .Y(n7843) );
  CLKBUFX3 U11576 ( .A(n7865), .Y(n7863) );
  CLKBUFX3 U11577 ( .A(n7865), .Y(n7864) );
  CLKBUFX3 U11578 ( .A(n7985), .Y(n7986) );
  CLKBUFX3 U11579 ( .A(n8049), .Y(n8050) );
  CLKBUFX3 U11580 ( .A(n8061), .Y(n8062) );
  CLKBUFX3 U11581 ( .A(n8100), .Y(n8101) );
  CLKBUFX3 U11582 ( .A(n8113), .Y(n8114) );
  CLKBUFX3 U11583 ( .A(n8126), .Y(n8127) );
  CLKBUFX3 U11584 ( .A(n8138), .Y(n8139) );
  CLKBUFX3 U11585 ( .A(n7972), .Y(n7973) );
  CLKBUFX3 U11586 ( .A(n7807), .Y(n7826) );
  CLKBUFX3 U11587 ( .A(n3678), .Y(n7928) );
  CLKBUFX3 U11588 ( .A(n3691), .Y(n7825) );
  CLKBUFX3 U11589 ( .A(n7807), .Y(n7824) );
  CLKBUFX3 U11590 ( .A(n7928), .Y(n7927) );
  CLKBUFX3 U11591 ( .A(n7807), .Y(n7823) );
  CLKBUFX3 U11592 ( .A(n3678), .Y(n7926) );
  CLKBUFX3 U11593 ( .A(n7889), .Y(n7908) );
  CLKINVX1 U11594 ( .A(n7846), .Y(n7832) );
  CLKINVX1 U11595 ( .A(n7847), .Y(n7851) );
  CLKBUFX3 U11596 ( .A(n7699), .Y(n7698) );
  CLKBUFX3 U11597 ( .A(n7689), .Y(n7688) );
  CLKBUFX3 U11598 ( .A(n7693), .Y(n7692) );
  CLKBUFX3 U11599 ( .A(n7695), .Y(n7694) );
  CLKBUFX3 U11600 ( .A(n7669), .Y(n7668) );
  CLKBUFX3 U11601 ( .A(n7671), .Y(n7670) );
  CLKBUFX3 U11602 ( .A(n7673), .Y(n7672) );
  CLKBUFX3 U11603 ( .A(n7677), .Y(n7676) );
  CLKBUFX3 U11604 ( .A(n7681), .Y(n7680) );
  CLKBUFX3 U11605 ( .A(n7683), .Y(n7682) );
  CLKBUFX3 U11606 ( .A(n7685), .Y(n7684) );
  CLKBUFX3 U11607 ( .A(n7697), .Y(n7696) );
  CLKBUFX3 U11608 ( .A(n6617), .Y(n7995) );
  CLKBUFX3 U11609 ( .A(n6618), .Y(n8007) );
  CLKBUFX3 U11610 ( .A(n8020), .Y(n8021) );
  CLKBUFX3 U11611 ( .A(n8033), .Y(n8034) );
  CLKBUFX3 U11612 ( .A(n8071), .Y(n8072) );
  CLKBUFX3 U11613 ( .A(n6619), .Y(n8084) );
  CLKBUFX3 U11614 ( .A(n6615), .Y(n8148) );
  CLKBUFX3 U11615 ( .A(n7995), .Y(n7996) );
  CLKBUFX3 U11616 ( .A(n8007), .Y(n8008) );
  CLKBUFX3 U11617 ( .A(n8084), .Y(n8085) );
  CLKBUFX3 U11618 ( .A(n8148), .Y(n8149) );
  CLKBUFX3 U11619 ( .A(n7995), .Y(n7997) );
  CLKBUFX3 U11620 ( .A(n8007), .Y(n8009) );
  CLKBUFX3 U11621 ( .A(n8021), .Y(n8022) );
  CLKBUFX3 U11622 ( .A(n8034), .Y(n8035) );
  CLKBUFX3 U11623 ( .A(n8072), .Y(n8073) );
  CLKBUFX3 U11624 ( .A(n8084), .Y(n8086) );
  CLKBUFX3 U11625 ( .A(n8148), .Y(n8150) );
  CLKBUFX3 U11626 ( .A(n8161), .Y(n8163) );
  CLKBUFX3 U11627 ( .A(n8061), .Y(n8063) );
  CLKBUFX3 U11628 ( .A(n8100), .Y(n8102) );
  CLKBUFX3 U11629 ( .A(n8113), .Y(n8115) );
  CLKBUFX3 U11630 ( .A(n8126), .Y(n8128) );
  CLKBUFX3 U11631 ( .A(n8138), .Y(n8140) );
  CLKBUFX3 U11632 ( .A(n7972), .Y(n7974) );
  CLKBUFX3 U11633 ( .A(n7650), .Y(n7635) );
  CLKBUFX3 U11634 ( .A(n7650), .Y(n7634) );
  CLKBUFX3 U11635 ( .A(n7650), .Y(n7633) );
  CLKBUFX3 U11636 ( .A(n7666), .Y(n7632) );
  CLKBUFX3 U11637 ( .A(n7666), .Y(n7631) );
  CLKBUFX3 U11638 ( .A(n7654), .Y(n7630) );
  CLKBUFX3 U11639 ( .A(n7651), .Y(n7629) );
  CLKBUFX3 U11640 ( .A(n7651), .Y(n7628) );
  CLKBUFX3 U11641 ( .A(n7651), .Y(n7627) );
  CLKBUFX3 U11642 ( .A(n7652), .Y(n7626) );
  CLKBUFX3 U11643 ( .A(n7652), .Y(n7625) );
  CLKBUFX3 U11644 ( .A(n7652), .Y(n7624) );
  CLKBUFX3 U11645 ( .A(n7665), .Y(n7623) );
  CLKBUFX3 U11646 ( .A(n7665), .Y(n7622) );
  CLKBUFX3 U11647 ( .A(n7663), .Y(n7621) );
  CLKBUFX3 U11648 ( .A(n7653), .Y(n7620) );
  CLKBUFX3 U11649 ( .A(n7653), .Y(n7619) );
  CLKBUFX3 U11650 ( .A(n7653), .Y(n7618) );
  CLKBUFX3 U11651 ( .A(n7654), .Y(n7617) );
  CLKBUFX3 U11652 ( .A(n7654), .Y(n7616) );
  CLKBUFX3 U11653 ( .A(n7654), .Y(n7615) );
  CLKBUFX3 U11654 ( .A(n7664), .Y(n7614) );
  CLKBUFX3 U11655 ( .A(n7569), .Y(n7613) );
  CLKBUFX3 U11656 ( .A(n8830), .Y(n7612) );
  CLKBUFX3 U11657 ( .A(n7655), .Y(n7611) );
  CLKBUFX3 U11658 ( .A(n7655), .Y(n7610) );
  CLKBUFX3 U11659 ( .A(n7655), .Y(n7609) );
  CLKBUFX3 U11660 ( .A(n7664), .Y(n7608) );
  CLKBUFX3 U11661 ( .A(n7664), .Y(n7607) );
  CLKBUFX3 U11662 ( .A(n7649), .Y(n7606) );
  CLKBUFX3 U11663 ( .A(n7656), .Y(n7605) );
  CLKBUFX3 U11664 ( .A(n7656), .Y(n7604) );
  CLKBUFX3 U11665 ( .A(n7656), .Y(n7603) );
  CLKBUFX3 U11666 ( .A(n7657), .Y(n7602) );
  CLKBUFX3 U11667 ( .A(n7657), .Y(n7601) );
  CLKBUFX3 U11668 ( .A(n7657), .Y(n7600) );
  CLKBUFX3 U11669 ( .A(n7663), .Y(n7599) );
  CLKBUFX3 U11670 ( .A(n7664), .Y(n7598) );
  CLKBUFX3 U11671 ( .A(n7655), .Y(n7597) );
  CLKBUFX3 U11672 ( .A(n7658), .Y(n7596) );
  CLKBUFX3 U11673 ( .A(n7658), .Y(n7595) );
  CLKBUFX3 U11674 ( .A(n7658), .Y(n7594) );
  CLKBUFX3 U11675 ( .A(n7659), .Y(n7593) );
  CLKBUFX3 U11676 ( .A(n7659), .Y(n7592) );
  CLKBUFX3 U11677 ( .A(n7659), .Y(n7591) );
  CLKBUFX3 U11678 ( .A(n7662), .Y(n7590) );
  CLKBUFX3 U11679 ( .A(n7662), .Y(n7589) );
  CLKBUFX3 U11680 ( .A(n7648), .Y(n7588) );
  CLKBUFX3 U11681 ( .A(n7661), .Y(n7587) );
  CLKBUFX3 U11682 ( .A(n7658), .Y(n7586) );
  CLKBUFX3 U11683 ( .A(n7659), .Y(n7585) );
  CLKBUFX3 U11684 ( .A(n7661), .Y(n7584) );
  CLKBUFX3 U11685 ( .A(n7661), .Y(n7583) );
  CLKBUFX3 U11686 ( .A(n7653), .Y(n7582) );
  CLKBUFX3 U11687 ( .A(n7661), .Y(n7581) );
  CLKBUFX3 U11688 ( .A(n7661), .Y(n7580) );
  CLKBUFX3 U11689 ( .A(n7567), .Y(n7579) );
  CLKBUFX3 U11690 ( .A(n7660), .Y(n7578) );
  CLKBUFX3 U11691 ( .A(n7651), .Y(n7577) );
  CLKBUFX3 U11692 ( .A(n7652), .Y(n7576) );
  CLKBUFX3 U11693 ( .A(n7660), .Y(n7575) );
  CLKBUFX3 U11694 ( .A(n7660), .Y(n7574) );
  CLKBUFX3 U11695 ( .A(n7567), .Y(n7573) );
  CLKBUFX3 U11696 ( .A(n7660), .Y(n7572) );
  CLKBUFX3 U11697 ( .A(n7656), .Y(n7571) );
  CLKBUFX3 U11698 ( .A(n7657), .Y(n7570) );
  CLKBUFX3 U11699 ( .A(n7648), .Y(n7641) );
  CLKBUFX3 U11700 ( .A(n7648), .Y(n7640) );
  CLKBUFX3 U11701 ( .A(n7648), .Y(n7639) );
  CLKBUFX3 U11702 ( .A(n7649), .Y(n7638) );
  CLKBUFX3 U11703 ( .A(n7649), .Y(n7637) );
  CLKBUFX3 U11704 ( .A(n7649), .Y(n7636) );
  CLKBUFX3 U11705 ( .A(n8335), .Y(n8325) );
  CLKBUFX3 U11706 ( .A(n8250), .Y(n8248) );
  CLKBUFX3 U11707 ( .A(n8303), .Y(n8301) );
  CLKBUFX3 U11708 ( .A(n8251), .Y(n8244) );
  CLKBUFX3 U11709 ( .A(n8251), .Y(n8245) );
  CLKBUFX3 U11710 ( .A(n8305), .Y(n8299) );
  CLKBUFX3 U11711 ( .A(n8250), .Y(n8247) );
  CLKBUFX3 U11712 ( .A(n8221), .Y(n8219) );
  CLKBUFX3 U11713 ( .A(n8222), .Y(n8216) );
  CLKBUFX3 U11714 ( .A(n8220), .Y(n8201) );
  CLKBUFX3 U11715 ( .A(n8221), .Y(n8220) );
  CLKBUFX3 U11716 ( .A(n8334), .Y(n8328) );
  CLKBUFX3 U11717 ( .A(n8335), .Y(n8326) );
  CLKBUFX3 U11718 ( .A(n8250), .Y(n8246) );
  CLKBUFX3 U11719 ( .A(n8304), .Y(n8300) );
  INVX3 U11720 ( .A(n8351), .Y(n8340) );
  INVX3 U11721 ( .A(n8351), .Y(n8347) );
  INVX3 U11722 ( .A(n8352), .Y(n8350) );
  CLKBUFX3 U11723 ( .A(n8215), .Y(n8211) );
  CLKBUFX3 U11724 ( .A(n8334), .Y(n8327) );
  CLKBUFX3 U11725 ( .A(n8333), .Y(n8330) );
  INVX3 U11726 ( .A(n8352), .Y(n8341) );
  CLKBUFX3 U11727 ( .A(n8222), .Y(n8217) );
  INVX3 U11728 ( .A(n8352), .Y(n8337) );
  CLKBUFX3 U11729 ( .A(n8250), .Y(n8249) );
  CLKBUFX3 U11730 ( .A(n8336), .Y(n8324) );
  CLKBUFX3 U11731 ( .A(n8333), .Y(n8331) );
  CLKBUFX3 U11732 ( .A(n8214), .Y(n8213) );
  CLKBUFX3 U11733 ( .A(n8334), .Y(n8329) );
  CLKBUFX3 U11734 ( .A(n8769), .Y(n7503) );
  CLKINVX1 U11735 ( .A(N25661), .Y(n8769) );
  CLKBUFX3 U11736 ( .A(n6981), .Y(n6982) );
  CLKBUFX3 U11737 ( .A(n7204), .Y(n7206) );
  CLKBUFX3 U11738 ( .A(n6981), .Y(n6983) );
  CLKBUFX3 U11739 ( .A(n6996), .Y(n6998) );
  CLKBUFX3 U11740 ( .A(n6996), .Y(n6997) );
  CLKBUFX3 U11741 ( .A(n6980), .Y(n6984) );
  INVX3 U11742 ( .A(n8351), .Y(n8339) );
  CLKBUFX3 U11743 ( .A(n6995), .Y(n6999) );
  INVX3 U11744 ( .A(n8352), .Y(n8342) );
  CLKBUFX3 U11745 ( .A(n6980), .Y(n6985) );
  CLKBUFX3 U11746 ( .A(n7203), .Y(n7208) );
  CLKBUFX3 U11747 ( .A(n6978), .Y(n6979) );
  CLKBUFX3 U11748 ( .A(n6992), .Y(n6994) );
  CLKBUFX3 U11749 ( .A(n6992), .Y(n6993) );
  INVX3 U11750 ( .A(n8352), .Y(n8338) );
  NAND2X1 U11751 ( .A(n3636), .B(n3637), .Y(n3572) );
  NAND2X1 U11752 ( .A(n2935), .B(n2936), .Y(n2808) );
  CLKBUFX3 U11753 ( .A(n8003), .Y(n8001) );
  CLKBUFX3 U11754 ( .A(n6585), .Y(n8003) );
  CLKBUFX3 U11755 ( .A(n8041), .Y(n8039) );
  CLKBUFX3 U11756 ( .A(n6576), .Y(n8041) );
  CLKBUFX3 U11757 ( .A(n8156), .Y(n8154) );
  CLKBUFX3 U11758 ( .A(n6586), .Y(n8156) );
  CLKBUFX3 U11759 ( .A(n6588), .Y(n8169) );
  CLKBUFX3 U11760 ( .A(n8046), .Y(n8045) );
  CLKBUFX3 U11761 ( .A(n8097), .Y(n8096) );
  CLKBUFX3 U11762 ( .A(n6584), .Y(n7988) );
  CLKBUFX3 U11763 ( .A(n6583), .Y(n8052) );
  CLKBUFX3 U11764 ( .A(n6607), .Y(n8064) );
  CLKBUFX3 U11765 ( .A(n6605), .Y(n8103) );
  CLKBUFX3 U11766 ( .A(n6606), .Y(n8116) );
  CLKBUFX3 U11767 ( .A(n6608), .Y(n8141) );
  NOR2BX1 U11768 ( .AN(n3636), .B(n3637), .Y(n3571) );
  NOR2BX1 U11769 ( .AN(n2935), .B(n2936), .Y(n2806) );
  CLKBUFX3 U11770 ( .A(n3153), .Y(n8058) );
  NOR2BX1 U11771 ( .AN(n3218), .B(n3219), .Y(n3153) );
  NOR2BX1 U11772 ( .AN(n2728), .B(n2729), .Y(n2599) );
  CLKBUFX3 U11773 ( .A(n3652), .Y(n7971) );
  CLKBUFX3 U11774 ( .A(n7975), .Y(n7976) );
  CLKBUFX3 U11775 ( .A(n7976), .Y(n7977) );
  CLKBUFX3 U11776 ( .A(n8104), .Y(n8105) );
  CLKBUFX3 U11777 ( .A(n8130), .Y(n8131) );
  CLKBUFX3 U11778 ( .A(n8027), .Y(n8028) );
  NOR2X1 U11779 ( .A(n8850), .B(n8849), .Y(n4844) );
  NAND2X1 U11780 ( .A(n4859), .B(n8849), .Y(n3498) );
  NAND2X1 U11781 ( .A(n8846), .B(n2936), .Y(n3671) );
  NAND3X1 U11782 ( .A(n8852), .B(n8851), .C(n4844), .Y(n4853) );
  CLKINVX1 U11783 ( .A(n4848), .Y(n8846) );
  CLKINVX1 U11784 ( .A(n4860), .Y(n8847) );
  CLKBUFX3 U11785 ( .A(n8080), .Y(n8083) );
  CLKBUFX3 U11786 ( .A(n3080), .Y(n8080) );
  CLKBUFX3 U11787 ( .A(n7867), .Y(n7886) );
  CLKBUFX3 U11788 ( .A(n3676), .Y(n7929) );
  CLKBUFX3 U11789 ( .A(n3695), .Y(n7767) );
  CLKBUFX3 U11790 ( .A(n6582), .Y(n7991) );
  NAND2X1 U11791 ( .A(n3639), .B(n3637), .Y(n3663) );
  CLKBUFX3 U11792 ( .A(n8860), .Y(n7761) );
  CLKBUFX3 U11793 ( .A(n8860), .Y(n7762) );
  CLKBUFX3 U11794 ( .A(n8860), .Y(n7763) );
  CLKBUFX3 U11795 ( .A(n8067), .Y(n8070) );
  CLKBUFX3 U11796 ( .A(n3149), .Y(n8067) );
  CLKBUFX3 U11797 ( .A(n6602), .Y(n8019) );
  CLKBUFX3 U11798 ( .A(n7784), .Y(n7805) );
  CLKBUFX3 U11799 ( .A(n7867), .Y(n7887) );
  CLKBUFX3 U11800 ( .A(n7783), .Y(n7804) );
  CLKBUFX3 U11801 ( .A(n8333), .Y(n8332) );
  CLKBUFX3 U11802 ( .A(n6611), .Y(n8029) );
  CLKBUFX3 U11803 ( .A(n6610), .Y(n8157) );
  CLKBUFX3 U11804 ( .A(n3667), .Y(n7944) );
  NOR2BX1 U11805 ( .AN(n2731), .B(n7700), .Y(n3667) );
  CLKBUFX3 U11806 ( .A(n3659), .Y(n7962) );
  NOR2BX1 U11807 ( .AN(n3293), .B(n8858), .Y(n3659) );
  NOR2BX1 U11808 ( .AN(n3221), .B(n8855), .Y(n3660) );
  CLKBUFX3 U11809 ( .A(n7784), .Y(n7806) );
  CLKBUFX3 U11810 ( .A(n7867), .Y(n7888) );
  CLKBUFX3 U11811 ( .A(n7374), .Y(n7367) );
  CLKBUFX3 U11812 ( .A(n7374), .Y(n7368) );
  CLKBUFX3 U11813 ( .A(n7374), .Y(n7369) );
  CLKBUFX3 U11814 ( .A(n7374), .Y(n7370) );
  CLKBUFX3 U11815 ( .A(n7374), .Y(n7371) );
  CLKBUFX3 U11816 ( .A(n7374), .Y(n7372) );
  CLKBUFX3 U11817 ( .A(n7374), .Y(n7373) );
  CLKBUFX3 U11818 ( .A(outCount_next[3]), .Y(n7357) );
  CLKINVX1 U11819 ( .A(n3219), .Y(n8855) );
  CLKBUFX3 U11820 ( .A(n215), .Y(n8376) );
  CLKBUFX3 U11821 ( .A(n215), .Y(n8375) );
  CLKBUFX3 U11822 ( .A(n218), .Y(n8374) );
  CLKBUFX3 U11823 ( .A(n218), .Y(n8373) );
  CLKBUFX3 U11824 ( .A(n222), .Y(n8372) );
  CLKBUFX3 U11825 ( .A(n222), .Y(n8371) );
  CLKBUFX3 U11826 ( .A(n226), .Y(n8370) );
  CLKBUFX3 U11827 ( .A(n226), .Y(n8369) );
  CLKBUFX3 U11828 ( .A(n230), .Y(n8368) );
  CLKBUFX3 U11829 ( .A(n230), .Y(n8367) );
  CLKBUFX3 U11830 ( .A(n234), .Y(n8366) );
  CLKBUFX3 U11831 ( .A(n234), .Y(n8365) );
  CLKBUFX3 U11832 ( .A(n164), .Y(n8394) );
  CLKBUFX3 U11833 ( .A(n164), .Y(n8393) );
  CLKBUFX3 U11834 ( .A(n183), .Y(n8392) );
  CLKBUFX3 U11835 ( .A(n183), .Y(n8391) );
  CLKBUFX3 U11836 ( .A(n187), .Y(n8390) );
  CLKBUFX3 U11837 ( .A(n187), .Y(n8389) );
  CLKBUFX3 U11838 ( .A(n191), .Y(n8388) );
  CLKBUFX3 U11839 ( .A(n191), .Y(n8387) );
  CLKBUFX3 U11840 ( .A(n195), .Y(n8386) );
  CLKBUFX3 U11841 ( .A(n195), .Y(n8385) );
  CLKBUFX3 U11842 ( .A(n199), .Y(n8384) );
  CLKBUFX3 U11843 ( .A(n199), .Y(n8383) );
  CLKBUFX3 U11844 ( .A(n203), .Y(n8382) );
  CLKBUFX3 U11845 ( .A(n203), .Y(n8381) );
  CLKBUFX3 U11846 ( .A(n207), .Y(n8380) );
  CLKBUFX3 U11847 ( .A(n207), .Y(n8379) );
  CLKBUFX3 U11848 ( .A(n211), .Y(n8378) );
  CLKBUFX3 U11849 ( .A(n211), .Y(n8377) );
  CLKBUFX3 U11850 ( .A(n238), .Y(n8364) );
  CLKBUFX3 U11851 ( .A(n238), .Y(n8363) );
  CLKBUFX3 U11852 ( .A(n7827), .Y(n7833) );
  CLKBUFX3 U11853 ( .A(n7847), .Y(n7852) );
  CLKBUFX3 U11854 ( .A(n7827), .Y(n7834) );
  CLKBUFX3 U11855 ( .A(n7847), .Y(n7853) );
  CLKBUFX3 U11856 ( .A(outCount_next[2]), .Y(n7359) );
  CLKBUFX3 U11857 ( .A(outCount_next[2]), .Y(n7360) );
  CLKBUFX3 U11858 ( .A(n3691), .Y(n7807) );
  CLKBUFX3 U11859 ( .A(n3680), .Y(n7889) );
  CLKBUFX3 U11860 ( .A(n3689), .Y(n7846) );
  CLKBUFX3 U11861 ( .A(n3687), .Y(n7866) );
  CLKBUFX3 U11862 ( .A(n7827), .Y(n7845) );
  CLKBUFX3 U11863 ( .A(n7827), .Y(n7844) );
  CLKBUFX3 U11864 ( .A(n7847), .Y(n7865) );
  CLKBUFX3 U11865 ( .A(n6720), .Y(n7686) );
  CLKBUFX3 U11866 ( .A(n6722), .Y(n7690) );
  CLKBUFX3 U11867 ( .A(n6727), .Y(n7674) );
  CLKBUFX3 U11868 ( .A(n6729), .Y(n7678) );
  CLKBUFX3 U11869 ( .A(n6591), .Y(n7985) );
  CLKBUFX3 U11870 ( .A(n6592), .Y(n8049) );
  CLKBUFX3 U11871 ( .A(n6593), .Y(n8061) );
  CLKBUFX3 U11872 ( .A(n6599), .Y(n8100) );
  CLKBUFX3 U11873 ( .A(n6598), .Y(n8113) );
  CLKBUFX3 U11874 ( .A(n6600), .Y(n8126) );
  CLKBUFX3 U11875 ( .A(n6594), .Y(n8138) );
  CLKBUFX3 U11876 ( .A(n6596), .Y(n7972) );
  CLKBUFX3 U11877 ( .A(n6612), .Y(n8020) );
  CLKBUFX3 U11878 ( .A(n6613), .Y(n8033) );
  CLKBUFX3 U11879 ( .A(n6614), .Y(n8071) );
  CLKBUFX3 U11880 ( .A(n6616), .Y(n8161) );
  CLKBUFX3 U11881 ( .A(n8401), .Y(n8400) );
  NOR2BX1 U11882 ( .AN(N34877), .B(n8401), .Y(xCount_next[0]) );
  CLKBUFX3 U11883 ( .A(n7985), .Y(n7987) );
  CLKBUFX3 U11884 ( .A(n8049), .Y(n8051) );
  CLKBUFX3 U11885 ( .A(n7569), .Y(n7646) );
  CLKBUFX3 U11886 ( .A(n7569), .Y(n7645) );
  CLKBUFX3 U11887 ( .A(n7568), .Y(n7644) );
  CLKBUFX3 U11888 ( .A(n7568), .Y(n7643) );
  CLKBUFX3 U11889 ( .A(n7650), .Y(n7642) );
  CLKBUFX3 U11890 ( .A(n7667), .Y(n7647) );
  CLKBUFX3 U11891 ( .A(n7667), .Y(n7650) );
  CLKBUFX3 U11892 ( .A(n7666), .Y(n7651) );
  CLKBUFX3 U11893 ( .A(n7666), .Y(n7652) );
  CLKBUFX3 U11894 ( .A(n7665), .Y(n7653) );
  CLKBUFX3 U11895 ( .A(n7665), .Y(n7654) );
  CLKBUFX3 U11896 ( .A(n7664), .Y(n7655) );
  CLKBUFX3 U11897 ( .A(n7663), .Y(n7656) );
  CLKBUFX3 U11898 ( .A(n7663), .Y(n7657) );
  CLKBUFX3 U11899 ( .A(n7662), .Y(n7658) );
  CLKBUFX3 U11900 ( .A(n7662), .Y(n7659) );
  CLKBUFX3 U11901 ( .A(n7667), .Y(n7648) );
  CLKBUFX3 U11902 ( .A(n7667), .Y(n7649) );
  CLKBUFX3 U11903 ( .A(n777), .Y(n8252) );
  CLKBUFX3 U11904 ( .A(n6711), .Y(n7710) );
  CLKBUFX3 U11905 ( .A(n6711), .Y(n7708) );
  CLKBUFX3 U11906 ( .A(n6711), .Y(n7707) );
  CLKBUFX3 U11907 ( .A(n6711), .Y(n7709) );
  CLKBUFX3 U11908 ( .A(n8223), .Y(n8215) );
  CLKBUFX3 U11909 ( .A(n6735), .Y(n8351) );
  CLKBUFX3 U11910 ( .A(n8859), .Y(n7750) );
  CLKBUFX3 U11911 ( .A(n262), .Y(n8357) );
  CLKBUFX3 U11912 ( .A(n8354), .Y(n8355) );
  CLKBUFX3 U11913 ( .A(n6597), .Y(n8354) );
  CLKBUFX3 U11914 ( .A(n6711), .Y(n7711) );
  CLKBUFX3 U11915 ( .A(n8223), .Y(n8214) );
  CLKBUFX3 U11916 ( .A(n7200), .Y(n7204) );
  CLKBUFX3 U11917 ( .A(n7212), .Y(n7216) );
  CLKBUFX3 U11918 ( .A(n6977), .Y(n6981) );
  CLKBUFX3 U11919 ( .A(n7226), .Y(n7224) );
  CLKBUFX3 U11920 ( .A(n7006), .Y(n7005) );
  CLKBUFX3 U11921 ( .A(N1763), .Y(n7223) );
  CLKBUFX3 U11922 ( .A(n7004), .Y(n7003) );
  CLKBUFX3 U11923 ( .A(n6991), .Y(n6996) );
  CLKBUFX3 U11924 ( .A(n262), .Y(n8356) );
  CLKBUFX3 U11925 ( .A(n6977), .Y(n6980) );
  CLKBUFX3 U11926 ( .A(n6991), .Y(n6995) );
  CLKBUFX3 U11927 ( .A(n7200), .Y(n7203) );
  CLKBUFX3 U11928 ( .A(n7212), .Y(n7215) );
  CLKBUFX3 U11929 ( .A(n6990), .Y(n6978) );
  CLKBUFX3 U11930 ( .A(n7002), .Y(n6992) );
  CLKBUFX3 U11931 ( .A(n7211), .Y(n7201) );
  CLKBUFX3 U11932 ( .A(n7217), .Y(n7213) );
  CLKBUFX3 U11933 ( .A(n6597), .Y(n8353) );
  NAND2X1 U11934 ( .A(n4821), .B(n4822), .Y(n3654) );
  NAND2X1 U11935 ( .A(n3007), .B(n3008), .Y(n2943) );
  NAND2X1 U11936 ( .A(n2800), .B(n2801), .Y(n2736) );
  NAND2X1 U11937 ( .A(n3290), .B(n3291), .Y(n3226) );
  NOR4X1 U11938 ( .A(n4828), .B(n4829), .C(n3648), .D(n4830), .Y(n4827) );
  NAND4X1 U11939 ( .A(n8876), .B(n8875), .C(n8874), .D(n8873), .Y(n4830) );
  NAND4X1 U11940 ( .A(n8868), .B(n8867), .C(n8866), .D(n8865), .Y(n4829) );
  NAND4X1 U11941 ( .A(n8864), .B(n8863), .C(n8862), .D(n8861), .Y(n4828) );
  CLKBUFX3 U11942 ( .A(n3649), .Y(n7975) );
  NOR2BX1 U11943 ( .AN(n4821), .B(n4822), .Y(n3652) );
  NOR2BX1 U11944 ( .AN(n3007), .B(n3008), .Y(n2942) );
  NOR2BX1 U11945 ( .AN(n2800), .B(n2801), .Y(n2735) );
  NAND2BX1 U11946 ( .AN(n8006), .B(n7502), .Y(n3431) );
  NAND2BX1 U11947 ( .AN(n8019), .B(n7502), .Y(n3362) );
  NAND2BX1 U11948 ( .AN(n8070), .B(n7502), .Y(n3081) );
  NAND2BX1 U11949 ( .AN(n8083), .B(n7502), .Y(n3010) );
  NOR2BX1 U11950 ( .AN(n3290), .B(n3291), .Y(n3225) );
  NAND4X1 U11951 ( .A(n8872), .B(n8871), .C(n8870), .D(n8869), .Y(n3648) );
  NOR2X1 U11952 ( .A(n8401), .B(n8861), .Y(xCount_next[31]) );
  NOR4X1 U11953 ( .A(n6595), .B(n6601), .C(n8849), .D(n8852), .Y(n3293) );
  NAND2X1 U11954 ( .A(n8848), .B(n3008), .Y(n3669) );
  NAND2X1 U11955 ( .A(n8847), .B(n2801), .Y(n3676) );
  AND4X1 U11956 ( .A(n3637), .B(n7803), .C(n4822), .D(n4873), .Y(n3700) );
  NOR3X1 U11957 ( .A(n7700), .B(n7768), .C(n7868), .Y(n4873) );
  NAND3XL U11958 ( .A(n6595), .B(n4840), .C(n4844), .Y(n4833) );
  NAND4XL U11959 ( .A(n8852), .B(n8849), .C(n6601), .D(n6595), .Y(n4848) );
  NAND3XL U11960 ( .A(n8852), .B(n6595), .C(n4844), .Y(n4860) );
  NOR2X1 U11961 ( .A(n8401), .B(n8866), .Y(xCount_next[26]) );
  NOR2X1 U11962 ( .A(n8401), .B(n8867), .Y(xCount_next[25]) );
  NOR2X1 U11963 ( .A(n8399), .B(n8862), .Y(xCount_next[30]) );
  NOR2X1 U11964 ( .A(n8399), .B(n8863), .Y(xCount_next[29]) );
  NOR2X1 U11965 ( .A(n8400), .B(n8864), .Y(xCount_next[28]) );
  NOR2X1 U11966 ( .A(n8401), .B(n8865), .Y(xCount_next[27]) );
  CLKBUFX3 U11967 ( .A(n3682), .Y(n7867) );
  NOR3BXL U11968 ( .AN(n4844), .B(n6595), .C(n8852), .Y(n2595) );
  OAI2BB2XL U11969 ( .B0(n4822), .B1(n4833), .A0N(n7704), .A1N(n3639), .Y(
        n6717) );
  CLKINVX1 U11970 ( .A(n6717), .Y(n3665) );
  OAI2BB2XL U11971 ( .B0(n4860), .B1(n2801), .A0N(n7700), .A1N(n2731), .Y(
        n6718) );
  CLKINVX1 U11972 ( .A(n6718), .Y(n3675) );
  NOR4X1 U11973 ( .A(n4840), .B(n6595), .C(n6601), .D(n4843), .Y(n3639) );
  NOR4X1 U11974 ( .A(n6601), .B(n4843), .C(n8851), .D(n8852), .Y(n3221) );
  NOR4X1 U11975 ( .A(n6595), .B(n4843), .C(n8850), .D(n8852), .Y(n2731) );
  INVX1 U11976 ( .A(n6601), .Y(n8850) );
  INVX3 U11977 ( .A(n4840), .Y(n8852) );
  NAND2X1 U11978 ( .A(n4861), .B(n8332), .Y(n2729) );
  NOR2X1 U11979 ( .A(n8401), .B(n8869), .Y(xCount_next[23]) );
  NOR2X1 U11980 ( .A(n8400), .B(n8870), .Y(xCount_next[22]) );
  NOR2X1 U11981 ( .A(n8400), .B(n8872), .Y(xCount_next[20]) );
  NOR2X1 U11982 ( .A(n8400), .B(n8874), .Y(xCount_next[18]) );
  NOR2X1 U11983 ( .A(n135), .B(n8868), .Y(xCount_next[24]) );
  NOR2X1 U11984 ( .A(n8399), .B(n8871), .Y(xCount_next[21]) );
  NOR2X1 U11985 ( .A(n135), .B(n8873), .Y(xCount_next[19]) );
  CLKBUFX3 U11986 ( .A(n3693), .Y(n7784) );
  CLKBUFX3 U11987 ( .A(n3693), .Y(n7783) );
  NAND2X1 U11988 ( .A(n4854), .B(n8352), .Y(n2936) );
  NAND2X1 U11989 ( .A(n4854), .B(n8332), .Y(n3691) );
  NAND2X1 U11990 ( .A(n4849), .B(n8332), .Y(n3680) );
  CLKINVX1 U11991 ( .A(n3291), .Y(n8858) );
  CLKBUFX3 U11992 ( .A(N35192), .Y(n8403) );
  CLKBUFX3 U11993 ( .A(N35192), .Y(n8402) );
  AND2X2 U11994 ( .A(n3220), .B(n2524), .Y(n185) );
  AND2X2 U11995 ( .A(n2523), .B(n2524), .Y(n240) );
  NOR2X1 U11996 ( .A(n8400), .B(n8875), .Y(xCount_next[17]) );
  NOR2X1 U11997 ( .A(n8400), .B(n8876), .Y(xCount_next[16]) );
  NOR2X1 U11998 ( .A(n8400), .B(n8877), .Y(xCount_next[12]) );
  CLKBUFX3 U11999 ( .A(n7358), .Y(n7356) );
  CLKBUFX3 U12000 ( .A(outCount_next[3]), .Y(n7358) );
  CLKBUFX3 U12001 ( .A(n3689), .Y(n7827) );
  CLKBUFX3 U12002 ( .A(n3687), .Y(n7847) );
  CLKBUFX3 U12003 ( .A(n8399), .Y(n8401) );
  CLKBUFX3 U12004 ( .A(n135), .Y(n8399) );
  NOR2BX1 U12005 ( .AN(N34880), .B(n8401), .Y(xCount_next[3]) );
  NOR2BX1 U12006 ( .AN(N34879), .B(n8401), .Y(xCount_next[2]) );
  NOR2BX1 U12007 ( .AN(N34878), .B(n8401), .Y(xCount_next[1]) );
  NOR2X1 U12008 ( .A(n8399), .B(n8883), .Y(xCount_next[4]) );
  NOR2X1 U12009 ( .A(n135), .B(n8882), .Y(xCount_next[5]) );
  NOR2X1 U12010 ( .A(n8399), .B(n8878), .Y(xCount_next[11]) );
  NOR2X1 U12011 ( .A(n135), .B(n8879), .Y(xCount_next[10]) );
  NOR2X1 U12012 ( .A(n8399), .B(n8880), .Y(xCount_next[7]) );
  NOR2X1 U12013 ( .A(n135), .B(n8881), .Y(xCount_next[6]) );
  CLKBUFX3 U12014 ( .A(n7567), .Y(n7666) );
  CLKBUFX3 U12015 ( .A(n7569), .Y(n7665) );
  CLKBUFX3 U12016 ( .A(n7569), .Y(n7664) );
  CLKBUFX3 U12017 ( .A(n7568), .Y(n7663) );
  CLKBUFX3 U12018 ( .A(n7568), .Y(n7662) );
  CLKBUFX3 U12019 ( .A(n7567), .Y(n7661) );
  CLKBUFX3 U12020 ( .A(n7567), .Y(n7660) );
  CLKBUFX3 U12021 ( .A(n8830), .Y(n7667) );
  OAI222XL U12022 ( .A0(n8938), .A1(n7941), .B0(n8478), .B1(n7938), .C0(n7936), 
        .C1(n8937), .Y(n3801) );
  OAI222XL U12023 ( .A0(n7956), .A1(n8935), .B0(n8942), .B1(n7953), .C0(n8478), 
        .C1(n7950), .Y(n3799) );
  OAI222XL U12024 ( .A0(n8930), .A1(n7941), .B0(n8473), .B1(n7938), .C0(n7936), 
        .C1(n8929), .Y(n3783) );
  OAI222XL U12025 ( .A0(n7956), .A1(n8927), .B0(n8934), .B1(n7953), .C0(n8473), 
        .C1(n7952), .Y(n3781) );
  OAI222XL U12026 ( .A0(n8922), .A1(n7941), .B0(n8468), .B1(n7938), .C0(n7936), 
        .C1(n8921), .Y(n3765) );
  OAI222XL U12027 ( .A0(n7956), .A1(n8919), .B0(n8926), .B1(n7953), .C0(n8468), 
        .C1(n7950), .Y(n3763) );
  OAI222XL U12028 ( .A0(n8914), .A1(n7941), .B0(n8463), .B1(n7938), .C0(n7936), 
        .C1(n8913), .Y(n3747) );
  OAI222XL U12029 ( .A0(n7956), .A1(n8911), .B0(n8918), .B1(n7953), .C0(n8463), 
        .C1(n7952), .Y(n3745) );
  OAI222XL U12030 ( .A0(n8906), .A1(n7941), .B0(n8453), .B1(n7938), .C0(n7936), 
        .C1(n8905), .Y(n3729) );
  OAI222XL U12031 ( .A0(n7956), .A1(n8903), .B0(n8910), .B1(n7955), .C0(n8453), 
        .C1(n7952), .Y(n3727) );
  OAI222XL U12032 ( .A0(n8898), .A1(n7941), .B0(n8448), .B1(n7938), .C0(n7936), 
        .C1(n8897), .Y(n3711) );
  OAI222XL U12033 ( .A0(n7956), .A1(n8895), .B0(n8902), .B1(n7954), .C0(n8448), 
        .C1(n7950), .Y(n3709) );
  OAI222XL U12034 ( .A0(n8890), .A1(n7941), .B0(n8458), .B1(n7938), .C0(n7936), 
        .C1(n8889), .Y(n3668) );
  OAI222XL U12035 ( .A0(n7956), .A1(n8887), .B0(n8894), .B1(n7953), .C0(n8458), 
        .C1(n7952), .Y(n3661) );
  OAI222XL U12036 ( .A0(n7487), .A1(n8002), .B0(n3509), .B1(n7998), .C0(n7507), 
        .C1(n7997), .Y(N27993) );
  OAI222XL U12037 ( .A0(n7487), .A1(n8015), .B0(n3441), .B1(n8010), .C0(n7507), 
        .C1(n8009), .Y(N28057) );
  OAI222XL U12038 ( .A0(n7487), .A1(n8028), .B0(n3372), .B1(n8023), .C0(n7507), 
        .C1(n8022), .Y(N28121) );
  OAI222XL U12039 ( .A0(n7487), .A1(n8041), .B0(n3304), .B1(n8036), .C0(n7507), 
        .C1(n8035), .Y(N28185) );
  OAI222XL U12040 ( .A0(n7487), .A1(n8079), .B0(n3091), .B1(n8074), .C0(n7507), 
        .C1(n8073), .Y(N28377) );
  OAI222XL U12041 ( .A0(n7487), .A1(n8092), .B0(n3020), .B1(n8087), .C0(n7507), 
        .C1(n8086), .Y(N28441) );
  OAI222XL U12042 ( .A0(n7487), .A1(n8155), .B0(n2537), .B1(n8151), .C0(n7507), 
        .C1(n8150), .Y(N28761) );
  OAI222XL U12043 ( .A0(n7487), .A1(n8168), .B0(n8165), .B1(n2353), .C0(n8163), 
        .C1(n7507), .Y(N28825) );
  OAI222XL U12044 ( .A0(n7489), .A1(n8002), .B0(n3508), .B1(n7998), .C0(n7506), 
        .C1(n7997), .Y(N27994) );
  OAI222XL U12045 ( .A0(n7489), .A1(n8015), .B0(n3440), .B1(n8010), .C0(n7506), 
        .C1(n8009), .Y(N28058) );
  OAI222XL U12046 ( .A0(n7489), .A1(n8028), .B0(n3371), .B1(n8023), .C0(n7506), 
        .C1(n8022), .Y(N28122) );
  OAI222XL U12047 ( .A0(n7489), .A1(n8041), .B0(n3303), .B1(n8036), .C0(n7506), 
        .C1(n8035), .Y(N28186) );
  OAI222XL U12048 ( .A0(n7489), .A1(n8079), .B0(n3090), .B1(n8074), .C0(n7506), 
        .C1(n8073), .Y(N28378) );
  OAI222XL U12049 ( .A0(n7489), .A1(n8092), .B0(n3019), .B1(n8087), .C0(n7506), 
        .C1(n8086), .Y(N28442) );
  OAI222XL U12050 ( .A0(n7489), .A1(n8155), .B0(n2536), .B1(n8151), .C0(n7506), 
        .C1(n8150), .Y(N28762) );
  OAI222XL U12051 ( .A0(n7489), .A1(n8168), .B0(n8165), .B1(n2350), .C0(n8163), 
        .C1(n7506), .Y(N28826) );
  OAI222XL U12052 ( .A0(n7491), .A1(n8003), .B0(n3507), .B1(n7998), .C0(n7505), 
        .C1(n7996), .Y(N27995) );
  OAI222XL U12053 ( .A0(n7491), .A1(n8014), .B0(n3439), .B1(n8010), .C0(n7505), 
        .C1(n8008), .Y(N28059) );
  OAI222XL U12054 ( .A0(n7491), .A1(n8028), .B0(n3370), .B1(n8023), .C0(n7505), 
        .C1(n6612), .Y(N28123) );
  OAI222XL U12055 ( .A0(n7491), .A1(n8041), .B0(n3302), .B1(n8036), .C0(n7505), 
        .C1(n8035), .Y(N28187) );
  OAI222XL U12056 ( .A0(n7491), .A1(n8078), .B0(n3089), .B1(n8074), .C0(n7505), 
        .C1(n8071), .Y(N28379) );
  OAI222XL U12057 ( .A0(n7491), .A1(n3010), .B0(n3018), .B1(n8087), .C0(n7505), 
        .C1(n8085), .Y(N28443) );
  OAI222XL U12058 ( .A0(n7491), .A1(n8156), .B0(n2535), .B1(n8151), .C0(n7505), 
        .C1(n8149), .Y(N28763) );
  OAI222XL U12059 ( .A0(n7491), .A1(n8167), .B0(n8165), .B1(n2347), .C0(n8163), 
        .C1(n7505), .Y(N28827) );
  OAI222XL U12060 ( .A0(n7493), .A1(n8002), .B0(n3506), .B1(n7998), .C0(n7504), 
        .C1(n7997), .Y(N27996) );
  OAI222XL U12061 ( .A0(n7493), .A1(n8015), .B0(n3438), .B1(n8010), .C0(n7504), 
        .C1(n8009), .Y(N28060) );
  OAI222XL U12062 ( .A0(n7493), .A1(n8028), .B0(n3369), .B1(n8023), .C0(n7504), 
        .C1(n8022), .Y(N28124) );
  OAI222XL U12063 ( .A0(n7493), .A1(n6576), .B0(n3301), .B1(n8036), .C0(n7504), 
        .C1(n8035), .Y(N28188) );
  OAI222XL U12064 ( .A0(n7493), .A1(n8079), .B0(n3088), .B1(n8074), .C0(n7504), 
        .C1(n8073), .Y(N28380) );
  OAI222XL U12065 ( .A0(n7493), .A1(n8092), .B0(n3017), .B1(n8087), .C0(n7504), 
        .C1(n8086), .Y(N28444) );
  OAI222XL U12066 ( .A0(n7493), .A1(n8155), .B0(n2534), .B1(n8151), .C0(n7504), 
        .C1(n8150), .Y(N28764) );
  OAI222XL U12067 ( .A0(n7493), .A1(n8168), .B0(n8165), .B1(n2344), .C0(n8161), 
        .C1(n7504), .Y(N28828) );
  OAI222XL U12068 ( .A0(n7495), .A1(n8001), .B0(n3505), .B1(n7998), .C0(n7503), 
        .C1(n7995), .Y(N27997) );
  OAI222XL U12069 ( .A0(n7495), .A1(n8013), .B0(n3437), .B1(n8010), .C0(n7503), 
        .C1(n8007), .Y(N28061) );
  OAI222XL U12070 ( .A0(n7495), .A1(n8028), .B0(n3368), .B1(n8023), .C0(n7503), 
        .C1(n8021), .Y(N28125) );
  OAI222XL U12071 ( .A0(n7495), .A1(n8041), .B0(n3300), .B1(n8036), .C0(n7503), 
        .C1(n8034), .Y(N28189) );
  OAI222XL U12072 ( .A0(n7495), .A1(n8077), .B0(n3087), .B1(n8074), .C0(n7503), 
        .C1(n8072), .Y(N28381) );
  OAI222XL U12073 ( .A0(n7495), .A1(n8091), .B0(n3016), .B1(n8087), .C0(n7503), 
        .C1(n8084), .Y(N28445) );
  OAI222XL U12074 ( .A0(n7495), .A1(n8156), .B0(n2533), .B1(n8151), .C0(n7503), 
        .C1(n8148), .Y(N28765) );
  OAI222XL U12075 ( .A0(n7495), .A1(n8167), .B0(n8165), .B1(n2341), .C0(n8163), 
        .C1(n7503), .Y(N28829) );
  OAI222XL U12076 ( .A0(n7497), .A1(n8002), .B0(n3504), .B1(n7998), .C0(n7564), 
        .C1(n7995), .Y(N27998) );
  OAI222XL U12077 ( .A0(n7497), .A1(n8013), .B0(n3436), .B1(n8010), .C0(n7564), 
        .C1(n8007), .Y(N28062) );
  OAI222XL U12078 ( .A0(n7497), .A1(n8028), .B0(n3367), .B1(n8023), .C0(n7564), 
        .C1(n8021), .Y(N28126) );
  OAI222XL U12079 ( .A0(n7497), .A1(n6576), .B0(n3299), .B1(n8036), .C0(n7565), 
        .C1(n8034), .Y(N28190) );
  OAI222XL U12080 ( .A0(n7497), .A1(n8077), .B0(n3086), .B1(n8074), .C0(n7565), 
        .C1(n8072), .Y(N28382) );
  OAI222XL U12081 ( .A0(n7497), .A1(n8091), .B0(n3015), .B1(n8087), .C0(n7565), 
        .C1(n8084), .Y(N28446) );
  OAI222XL U12082 ( .A0(n7497), .A1(n8155), .B0(n2532), .B1(n8151), .C0(n7564), 
        .C1(n8148), .Y(N28766) );
  OAI222XL U12083 ( .A0(n7497), .A1(n8168), .B0(n8165), .B1(n2338), .C0(n8162), 
        .C1(n7564), .Y(N28830) );
  OAI222XL U12084 ( .A0(n7499), .A1(n8001), .B0(n3503), .B1(n7998), .C0(n7564), 
        .C1(n7995), .Y(N27999) );
  OAI222XL U12085 ( .A0(n7499), .A1(n8013), .B0(n3435), .B1(n8010), .C0(n7565), 
        .C1(n8007), .Y(N28063) );
  OAI222XL U12086 ( .A0(n7499), .A1(n8028), .B0(n3366), .B1(n8023), .C0(n7565), 
        .C1(n8021), .Y(N28127) );
  OAI222XL U12087 ( .A0(n7499), .A1(n6576), .B0(n3298), .B1(n8036), .C0(n7565), 
        .C1(n8034), .Y(N28191) );
  OAI222XL U12088 ( .A0(n7499), .A1(n8077), .B0(n3085), .B1(n8074), .C0(n7565), 
        .C1(n8072), .Y(N28383) );
  OAI222XL U12089 ( .A0(n7499), .A1(n8091), .B0(n3014), .B1(n8087), .C0(n7564), 
        .C1(n8084), .Y(N28447) );
  OAI222XL U12090 ( .A0(n7499), .A1(n8156), .B0(n2531), .B1(n8151), .C0(n7564), 
        .C1(n8148), .Y(N28767) );
  OAI222XL U12091 ( .A0(n7499), .A1(n8167), .B0(n8165), .B1(n2335), .C0(n8162), 
        .C1(n7564), .Y(N28831) );
  OAI222XL U12092 ( .A0(n7501), .A1(n8002), .B0(n3500), .B1(n7998), .C0(n7564), 
        .C1(n7995), .Y(N28000) );
  OAI222XL U12093 ( .A0(n7501), .A1(n8013), .B0(n3432), .B1(n8010), .C0(n7564), 
        .C1(n8007), .Y(N28064) );
  OAI222XL U12094 ( .A0(n7501), .A1(n8028), .B0(n3363), .B1(n8023), .C0(n7565), 
        .C1(n8021), .Y(N28128) );
  OAI222XL U12095 ( .A0(n7501), .A1(n8041), .B0(n3295), .B1(n8036), .C0(n7565), 
        .C1(n8034), .Y(N28192) );
  OAI222XL U12096 ( .A0(n7501), .A1(n8077), .B0(n3082), .B1(n8074), .C0(n7565), 
        .C1(n8072), .Y(N28384) );
  OAI222XL U12097 ( .A0(n7501), .A1(n8091), .B0(n3011), .B1(n8087), .C0(n7565), 
        .C1(n8084), .Y(N28448) );
  OAI222XL U12098 ( .A0(n7501), .A1(n8155), .B0(n2528), .B1(n8151), .C0(n7564), 
        .C1(n8148), .Y(N28768) );
  OAI222XL U12099 ( .A0(n7501), .A1(n8168), .B0(n8165), .B1(n2331), .C0(n8162), 
        .C1(n7564), .Y(N28832) );
  OAI222XL U12100 ( .A0(n8473), .A1(n7932), .B0(n7931), .B1(n8928), .C0(n8006), 
        .C1(n3439), .Y(n3786) );
  OAI222XL U12101 ( .A0(n8468), .A1(n7932), .B0(n7931), .B1(n8920), .C0(n8006), 
        .C1(n3438), .Y(n3768) );
  OAI222XL U12102 ( .A0(n8463), .A1(n7932), .B0(n7931), .B1(n8912), .C0(n8006), 
        .C1(n3437), .Y(n3750) );
  OAI222XL U12103 ( .A0(n8453), .A1(n7932), .B0(n7929), .B1(n8904), .C0(n8006), 
        .C1(n3436), .Y(n3732) );
  OAI222XL U12104 ( .A0(n8448), .A1(n7932), .B0(n7930), .B1(n8896), .C0(n8006), 
        .C1(n3435), .Y(n3714) );
  OAI222XL U12105 ( .A0(n8483), .A1(n7932), .B0(n7929), .B1(n8944), .C0(n8006), 
        .C1(n3441), .Y(n3822) );
  OAI222XL U12106 ( .A0(n8478), .A1(n7932), .B0(n7930), .B1(n8936), .C0(n8006), 
        .C1(n3440), .Y(n3804) );
  OAI222XL U12107 ( .A0(n8458), .A1(n7932), .B0(n7931), .B1(n8888), .C0(n3432), 
        .C1(n8004), .Y(n3674) );
  OAI221XL U12108 ( .A0(n7487), .A1(n7990), .B0(n7507), .B1(n7987), .C0(n3579), 
        .Y(N27929) );
  OAI221XL U12109 ( .A0(n7487), .A1(n8054), .B0(n7507), .B1(n8051), .C0(n3233), 
        .Y(N28249) );
  OAI221XL U12110 ( .A0(n7487), .A1(n8105), .B0(n7507), .B1(n6599), .C0(n2950), 
        .Y(N28505) );
  OAI221XL U12111 ( .A0(n7487), .A1(n8116), .B0(n7507), .B1(n6598), .C0(n2821), 
        .Y(N28569) );
  OAI221XL U12112 ( .A0(n7487), .A1(n8131), .B0(n7507), .B1(n6600), .C0(n2743), 
        .Y(N28633) );
  OAI221XL U12113 ( .A0(n7487), .A1(n7975), .B0(n7507), .B1(n7974), .C0(n3811), 
        .Y(N27865) );
  OAI221XL U12114 ( .A0(n7489), .A1(n7990), .B0(n7506), .B1(n7987), .C0(n3578), 
        .Y(N27930) );
  OAI221XL U12115 ( .A0(n7489), .A1(n8054), .B0(n7506), .B1(n8051), .C0(n3232), 
        .Y(N28250) );
  OAI221XL U12116 ( .A0(n7489), .A1(n8105), .B0(n7506), .B1(n6599), .C0(n2949), 
        .Y(N28506) );
  OAI221XL U12117 ( .A0(n7489), .A1(n8116), .B0(n7506), .B1(n6598), .C0(n2819), 
        .Y(N28570) );
  OAI221XL U12118 ( .A0(n7489), .A1(n8131), .B0(n7506), .B1(n6600), .C0(n2742), 
        .Y(N28634) );
  OAI221XL U12119 ( .A0(n7489), .A1(n7975), .B0(n7506), .B1(n7974), .C0(n3793), 
        .Y(N27866) );
  OAI221XL U12120 ( .A0(n7491), .A1(n7990), .B0(n7505), .B1(n7987), .C0(n3577), 
        .Y(N27931) );
  OAI221XL U12121 ( .A0(n7491), .A1(n8054), .B0(n7505), .B1(n8051), .C0(n3231), 
        .Y(N28251) );
  OAI221XL U12122 ( .A0(n7491), .A1(n8105), .B0(n7505), .B1(n8101), .C0(n2948), 
        .Y(N28507) );
  OAI221XL U12123 ( .A0(n7491), .A1(n8116), .B0(n7505), .B1(n8114), .C0(n2817), 
        .Y(N28571) );
  OAI221XL U12124 ( .A0(n7491), .A1(n8131), .B0(n7505), .B1(n8127), .C0(n2741), 
        .Y(N28635) );
  OAI221XL U12125 ( .A0(n7491), .A1(n7976), .B0(n7505), .B1(n7973), .C0(n3775), 
        .Y(N27867) );
  OAI221XL U12126 ( .A0(n7493), .A1(n7988), .B0(n7504), .B1(n7987), .C0(n3576), 
        .Y(N27932) );
  OAI221XL U12127 ( .A0(n7493), .A1(n8052), .B0(n7504), .B1(n8051), .C0(n3230), 
        .Y(N28252) );
  OAI221XL U12128 ( .A0(n7493), .A1(n8105), .B0(n7504), .B1(n6599), .C0(n2947), 
        .Y(N28508) );
  OAI221XL U12129 ( .A0(n7493), .A1(n8116), .B0(n7504), .B1(n6598), .C0(n2815), 
        .Y(N28572) );
  OAI221XL U12130 ( .A0(n7493), .A1(n8131), .B0(n7504), .B1(n8126), .C0(n2740), 
        .Y(N28636) );
  OAI221XL U12131 ( .A0(n7493), .A1(n7975), .B0(n7504), .B1(n7972), .C0(n3757), 
        .Y(N27868) );
  OAI221XL U12132 ( .A0(n7495), .A1(n7988), .B0(n7503), .B1(n7987), .C0(n3575), 
        .Y(N27933) );
  OAI221XL U12133 ( .A0(n7495), .A1(n8052), .B0(n7503), .B1(n8051), .C0(n3229), 
        .Y(N28253) );
  OAI221XL U12134 ( .A0(n7495), .A1(n8105), .B0(n7503), .B1(n8101), .C0(n2946), 
        .Y(N28509) );
  OAI221XL U12135 ( .A0(n7495), .A1(n8116), .B0(n7503), .B1(n8114), .C0(n2813), 
        .Y(N28573) );
  OAI221XL U12136 ( .A0(n7495), .A1(n8131), .B0(n7503), .B1(n8127), .C0(n2739), 
        .Y(N28637) );
  OAI221XL U12137 ( .A0(n7495), .A1(n7976), .B0(n7503), .B1(n6596), .C0(n3739), 
        .Y(N27869) );
  OAI221XL U12138 ( .A0(n7497), .A1(n7988), .B0(n7566), .B1(n7987), .C0(n3574), 
        .Y(N27934) );
  OAI221XL U12139 ( .A0(n7497), .A1(n8052), .B0(n7566), .B1(n8051), .C0(n3228), 
        .Y(N28254) );
  OAI221XL U12140 ( .A0(n7497), .A1(n8105), .B0(n7566), .B1(n8102), .C0(n2945), 
        .Y(N28510) );
  OAI221XL U12141 ( .A0(n7497), .A1(n8117), .B0(n7566), .B1(n8113), .C0(n2811), 
        .Y(N28574) );
  OAI221XL U12142 ( .A0(n7497), .A1(n8131), .B0(n7564), .B1(n8128), .C0(n2738), 
        .Y(N28638) );
  OAI221XL U12143 ( .A0(n7497), .A1(n7977), .B0(n7564), .B1(n6596), .C0(n3721), 
        .Y(N27870) );
  OAI221XL U12144 ( .A0(n7499), .A1(n7988), .B0(n7566), .B1(n7987), .C0(n3573), 
        .Y(N27935) );
  OAI221XL U12145 ( .A0(n7499), .A1(n8054), .B0(n7566), .B1(n8051), .C0(n3227), 
        .Y(N28255) );
  OAI221XL U12146 ( .A0(n7499), .A1(n8105), .B0(n7566), .B1(n8100), .C0(n2944), 
        .Y(N28511) );
  OAI221XL U12147 ( .A0(n7499), .A1(n8117), .B0(n7565), .B1(n8115), .C0(n2809), 
        .Y(N28575) );
  OAI221XL U12148 ( .A0(n7499), .A1(n8131), .B0(n8768), .B1(n8128), .C0(n2737), 
        .Y(N28639) );
  OAI221XL U12149 ( .A0(n7499), .A1(n7975), .B0(n7566), .B1(n6596), .C0(n3703), 
        .Y(N27871) );
  OAI221XL U12150 ( .A0(n7501), .A1(n7990), .B0(n7566), .B1(n7987), .C0(n3570), 
        .Y(N27936) );
  OAI221XL U12151 ( .A0(n7501), .A1(n8054), .B0(n7566), .B1(n8051), .C0(n3224), 
        .Y(N28256) );
  OAI221XL U12152 ( .A0(n7501), .A1(n8105), .B0(n7565), .B1(n8101), .C0(n2941), 
        .Y(N28512) );
  OAI221XL U12153 ( .A0(n7501), .A1(n8117), .B0(n7566), .B1(n8114), .C0(n2805), 
        .Y(N28576) );
  OAI221XL U12154 ( .A0(n7501), .A1(n8131), .B0(n8768), .B1(n8128), .C0(n2734), 
        .Y(N28640) );
  OAI221XL U12155 ( .A0(n7501), .A1(n7976), .B0(n7565), .B1(n6596), .C0(n3651), 
        .Y(N27872) );
  CLKBUFX3 U12156 ( .A(n268), .Y(n8307) );
  CLKBUFX3 U12157 ( .A(n786), .Y(n8182) );
  CLKBUFX3 U12158 ( .A(n779), .Y(n8224) );
  CLKBUFX3 U12159 ( .A(n775), .Y(n8278) );
  OAI222XL U12160 ( .A0(n8503), .A1(n7932), .B0(n7929), .B1(n8976), .C0(n8006), 
        .C1(n3445), .Y(n3894) );
  OAI222XL U12161 ( .A0(n7956), .A1(n8975), .B0(n8982), .B1(n7955), .C0(n8503), 
        .C1(n7952), .Y(n3889) );
  OAI222XL U12162 ( .A0(n8970), .A1(n7941), .B0(n8498), .B1(n7938), .C0(n7936), 
        .C1(n8969), .Y(n3873) );
  OAI222XL U12163 ( .A0(n7956), .A1(n8967), .B0(n8974), .B1(n7953), .C0(n8498), 
        .C1(n7952), .Y(n3871) );
  OAI222XL U12164 ( .A0(n8962), .A1(n7941), .B0(n8493), .B1(n7938), .C0(n7936), 
        .C1(n8961), .Y(n3855) );
  OAI222XL U12165 ( .A0(n7956), .A1(n8959), .B0(n8966), .B1(n7953), .C0(n8493), 
        .C1(n7950), .Y(n3853) );
  OAI222XL U12166 ( .A0(n8954), .A1(n7941), .B0(n8488), .B1(n7938), .C0(n7936), 
        .C1(n8953), .Y(n3837) );
  OAI222XL U12167 ( .A0(n7956), .A1(n8951), .B0(n8958), .B1(n7955), .C0(n8488), 
        .C1(n7952), .Y(n3835) );
  OAI222XL U12168 ( .A0(n8946), .A1(n7941), .B0(n8483), .B1(n7938), .C0(n7936), 
        .C1(n8945), .Y(n3819) );
  OAI222XL U12169 ( .A0(n7956), .A1(n8943), .B0(n8950), .B1(n7953), .C0(n8483), 
        .C1(n7950), .Y(n3817) );
  OAI222XL U12170 ( .A0(n7479), .A1(n8015), .B0(n3445), .B1(n8010), .C0(n7511), 
        .C1(n8009), .Y(N28053) );
  OAI222XL U12171 ( .A0(n7479), .A1(n8028), .B0(n3376), .B1(n8023), .C0(n7511), 
        .C1(n8022), .Y(N28117) );
  OAI222XL U12172 ( .A0(n7479), .A1(n8079), .B0(n3095), .B1(n8074), .C0(n7511), 
        .C1(n8073), .Y(N28373) );
  OAI222XL U12173 ( .A0(n7479), .A1(n8092), .B0(n3024), .B1(n8087), .C0(n7511), 
        .C1(n8086), .Y(N28437) );
  OAI222XL U12174 ( .A0(n7481), .A1(n8002), .B0(n3512), .B1(n7998), .C0(n7510), 
        .C1(n7997), .Y(N27990) );
  OAI222XL U12175 ( .A0(n7481), .A1(n8015), .B0(n3444), .B1(n8010), .C0(n7510), 
        .C1(n8009), .Y(N28054) );
  OAI222XL U12176 ( .A0(n7481), .A1(n3362), .B0(n3375), .B1(n8023), .C0(n7510), 
        .C1(n8022), .Y(N28118) );
  OAI222XL U12177 ( .A0(n7481), .A1(n8041), .B0(n3307), .B1(n8036), .C0(n7510), 
        .C1(n8035), .Y(N28182) );
  OAI222XL U12178 ( .A0(n7481), .A1(n8079), .B0(n3094), .B1(n8074), .C0(n7510), 
        .C1(n8073), .Y(N28374) );
  OAI222XL U12179 ( .A0(n7481), .A1(n8092), .B0(n3023), .B1(n8087), .C0(n7510), 
        .C1(n8086), .Y(N28438) );
  OAI222XL U12180 ( .A0(n7481), .A1(n8155), .B0(n2540), .B1(n8151), .C0(n7510), 
        .C1(n8150), .Y(N28758) );
  OAI222XL U12181 ( .A0(n7481), .A1(n8168), .B0(n8165), .B1(n2362), .C0(n8163), 
        .C1(n7510), .Y(N28822) );
  OAI222XL U12182 ( .A0(n7483), .A1(n8002), .B0(n3511), .B1(n7998), .C0(n7509), 
        .C1(n7997), .Y(N27991) );
  OAI222XL U12183 ( .A0(n7483), .A1(n8015), .B0(n3443), .B1(n8010), .C0(n7509), 
        .C1(n8009), .Y(N28055) );
  OAI222XL U12184 ( .A0(n7483), .A1(n8028), .B0(n3374), .B1(n8023), .C0(n7509), 
        .C1(n8022), .Y(N28119) );
  OAI222XL U12185 ( .A0(n7483), .A1(n8041), .B0(n3306), .B1(n8036), .C0(n7509), 
        .C1(n8035), .Y(N28183) );
  OAI222XL U12186 ( .A0(n7483), .A1(n8079), .B0(n3093), .B1(n8074), .C0(n7509), 
        .C1(n8073), .Y(N28375) );
  OAI222XL U12187 ( .A0(n7483), .A1(n8092), .B0(n3022), .B1(n8087), .C0(n7509), 
        .C1(n8086), .Y(N28439) );
  OAI222XL U12188 ( .A0(n7483), .A1(n8155), .B0(n2539), .B1(n8151), .C0(n7509), 
        .C1(n8150), .Y(N28759) );
  OAI222XL U12189 ( .A0(n7483), .A1(n8168), .B0(n8165), .B1(n2359), .C0(n8163), 
        .C1(n7509), .Y(N28823) );
  OAI222XL U12190 ( .A0(n7485), .A1(n8002), .B0(n3510), .B1(n7998), .C0(n7508), 
        .C1(n7997), .Y(N27992) );
  OAI222XL U12191 ( .A0(n7485), .A1(n8015), .B0(n3442), .B1(n8010), .C0(n7508), 
        .C1(n8009), .Y(N28056) );
  OAI222XL U12192 ( .A0(n7485), .A1(n8027), .B0(n3373), .B1(n8023), .C0(n7508), 
        .C1(n8022), .Y(N28120) );
  OAI222XL U12193 ( .A0(n7485), .A1(n8041), .B0(n3305), .B1(n8036), .C0(n7508), 
        .C1(n8035), .Y(N28184) );
  OAI222XL U12194 ( .A0(n7485), .A1(n8079), .B0(n3092), .B1(n8074), .C0(n7508), 
        .C1(n8073), .Y(N28376) );
  OAI222XL U12195 ( .A0(n7485), .A1(n8092), .B0(n3021), .B1(n8087), .C0(n7508), 
        .C1(n8086), .Y(N28440) );
  OAI222XL U12196 ( .A0(n7485), .A1(n8155), .B0(n2538), .B1(n8151), .C0(n7508), 
        .C1(n8150), .Y(N28760) );
  OAI222XL U12197 ( .A0(n7485), .A1(n8168), .B0(n8165), .B1(n2356), .C0(n8163), 
        .C1(n7508), .Y(N28824) );
  AOI221XL U12198 ( .A0(n8504), .A1(n8158), .B0(n8505), .B1(n8147), .C0(n3897), 
        .Y(n3885) );
  OAI222XL U12199 ( .A0(n8083), .A1(n3024), .B0(n8019), .B1(n3376), .C0(n8070), 
        .C1(n3095), .Y(n3897) );
  OAI222XL U12200 ( .A0(n8498), .A1(n7932), .B0(n7929), .B1(n8968), .C0(n8006), 
        .C1(n3444), .Y(n3876) );
  OAI222XL U12201 ( .A0(n8493), .A1(n7932), .B0(n7929), .B1(n8960), .C0(n8006), 
        .C1(n3443), .Y(n3858) );
  OAI222XL U12202 ( .A0(n8488), .A1(n7932), .B0(n3676), .B1(n8952), .C0(n8006), 
        .C1(n3442), .Y(n3840) );
  OAI221XL U12203 ( .A0(n7479), .A1(n7990), .B0(n7511), .B1(n7987), .C0(n3583), 
        .Y(N27925) );
  AOI2BB2X1 U12204 ( .B0(n7982), .B1(n7478), .A0N(n8982), .A1N(n7978), .Y(
        n3583) );
  OAI221XL U12205 ( .A0(n7479), .A1(n8054), .B0(n7511), .B1(n8051), .C0(n3237), 
        .Y(N28245) );
  AOI2BB2X1 U12206 ( .B0(n8046), .B1(n7478), .A0N(n8980), .A1N(n8042), .Y(
        n3237) );
  OAI221XL U12207 ( .A0(n7479), .A1(n8103), .B0(n7511), .B1(n8100), .C0(n2954), 
        .Y(N28501) );
  AOI2BB2X1 U12208 ( .B0(n8098), .B1(n7478), .A0N(n8978), .A1N(n8093), .Y(
        n2954) );
  OAI221XL U12209 ( .A0(n7479), .A1(n8116), .B0(n7511), .B1(n8113), .C0(n2829), 
        .Y(N28565) );
  AOI2BB2X1 U12210 ( .B0(n8111), .B1(n7478), .A0N(n8977), .A1N(n8106), .Y(
        n2829) );
  OAI221XL U12211 ( .A0(n7479), .A1(n6609), .B0(n7511), .B1(n8127), .C0(n2747), 
        .Y(N28629) );
  AOI2BB2X1 U12212 ( .B0(n8123), .B1(n7478), .A0N(n8976), .A1N(n8119), .Y(
        n2747) );
  OAI221XL U12213 ( .A0(n7479), .A1(n7975), .B0(n7511), .B1(n6596), .C0(n3883), 
        .Y(N27861) );
  AOI2BB2X1 U12214 ( .B0(n7970), .B1(n7478), .A0N(n8975), .A1N(n7966), .Y(
        n3883) );
  OAI221XL U12215 ( .A0(n7481), .A1(n7990), .B0(n7510), .B1(n7987), .C0(n3582), 
        .Y(N27926) );
  OAI221XL U12216 ( .A0(n7481), .A1(n8054), .B0(n7510), .B1(n8051), .C0(n3236), 
        .Y(N28246) );
  OAI221XL U12217 ( .A0(n7481), .A1(n8104), .B0(n7510), .B1(n8101), .C0(n2953), 
        .Y(N28502) );
  OAI221XL U12218 ( .A0(n7481), .A1(n8116), .B0(n7510), .B1(n8114), .C0(n2827), 
        .Y(N28566) );
  OAI221XL U12219 ( .A0(n7481), .A1(n8130), .B0(n7510), .B1(n8127), .C0(n2746), 
        .Y(N28630) );
  OAI221XL U12220 ( .A0(n7481), .A1(n7975), .B0(n7510), .B1(n6596), .C0(n3865), 
        .Y(N27862) );
  OAI221XL U12221 ( .A0(n7483), .A1(n7988), .B0(n7509), .B1(n7987), .C0(n3581), 
        .Y(N27927) );
  OAI221XL U12222 ( .A0(n7483), .A1(n8052), .B0(n7509), .B1(n8051), .C0(n3235), 
        .Y(N28247) );
  OAI221XL U12223 ( .A0(n7483), .A1(n8105), .B0(n7509), .B1(n8101), .C0(n2952), 
        .Y(N28503) );
  OAI221XL U12224 ( .A0(n7483), .A1(n8117), .B0(n7509), .B1(n8114), .C0(n2825), 
        .Y(N28567) );
  OAI221XL U12225 ( .A0(n7483), .A1(n8131), .B0(n7509), .B1(n8127), .C0(n2745), 
        .Y(N28631) );
  OAI221XL U12226 ( .A0(n7483), .A1(n7976), .B0(n7509), .B1(n7972), .C0(n3847), 
        .Y(N27863) );
  OAI221XL U12227 ( .A0(n7485), .A1(n7988), .B0(n7508), .B1(n7987), .C0(n3580), 
        .Y(N27928) );
  OAI221XL U12228 ( .A0(n7485), .A1(n8052), .B0(n7508), .B1(n8051), .C0(n3234), 
        .Y(N28248) );
  OAI221XL U12229 ( .A0(n7485), .A1(n8105), .B0(n7508), .B1(n8101), .C0(n2951), 
        .Y(N28504) );
  OAI221XL U12230 ( .A0(n7485), .A1(n8117), .B0(n7508), .B1(n8114), .C0(n2823), 
        .Y(N28568) );
  OAI221XL U12231 ( .A0(n7485), .A1(n8131), .B0(n7508), .B1(n8127), .C0(n2744), 
        .Y(N28632) );
  OAI221XL U12232 ( .A0(n7485), .A1(n7976), .B0(n7508), .B1(n7972), .C0(n3829), 
        .Y(N27864) );
  OA22X1 U12233 ( .A0(n7754), .A1(n968), .B0(n8340), .B1(n1542), .Y(n1541) );
  CLKBUFX3 U12234 ( .A(n268), .Y(n8306) );
  CLKBUFX3 U12235 ( .A(n6707), .Y(n8183) );
  OAI222XL U12236 ( .A0(n9002), .A1(n7942), .B0(n8518), .B1(n7939), .C0(n7935), 
        .C1(n9001), .Y(n3945) );
  OAI222XL U12237 ( .A0(n8994), .A1(n7942), .B0(n8513), .B1(n7939), .C0(n7935), 
        .C1(n8993), .Y(n3927) );
  OAI222XL U12238 ( .A0(n3662), .A1(n8991), .B0(n8998), .B1(n7955), .C0(n8513), 
        .C1(n7950), .Y(n3925) );
  OAI222XL U12239 ( .A0(n8508), .A1(n7933), .B0(n3676), .B1(n8984), .C0(n8006), 
        .C1(n3446), .Y(n3912) );
  OAI222XL U12240 ( .A0(n7956), .A1(n8983), .B0(n8990), .B1(n7954), .C0(n8508), 
        .C1(n7950), .Y(n3907) );
  OAI222XL U12241 ( .A0(n7473), .A1(n8002), .B0(n3516), .B1(n7999), .C0(n7514), 
        .C1(n7997), .Y(N27986) );
  OAI222XL U12242 ( .A0(n7473), .A1(n8015), .B0(n3448), .B1(n8010), .C0(n7514), 
        .C1(n8009), .Y(N28050) );
  OAI222XL U12243 ( .A0(n7473), .A1(n8027), .B0(n3379), .B1(n8023), .C0(n7514), 
        .C1(n8022), .Y(N28114) );
  OAI222XL U12244 ( .A0(n7473), .A1(n8041), .B0(n3311), .B1(n8037), .C0(n7514), 
        .C1(n8035), .Y(N28178) );
  OAI222XL U12245 ( .A0(n7473), .A1(n8079), .B0(n3098), .B1(n8075), .C0(n7514), 
        .C1(n8073), .Y(N28370) );
  OAI222XL U12246 ( .A0(n7473), .A1(n8092), .B0(n3027), .B1(n8088), .C0(n7514), 
        .C1(n8086), .Y(N28434) );
  OAI222XL U12247 ( .A0(n7473), .A1(n8155), .B0(n2544), .B1(n8152), .C0(n7514), 
        .C1(n8150), .Y(N28754) );
  OAI222XL U12248 ( .A0(n7473), .A1(n8168), .B0(n8164), .B1(n2374), .C0(n8163), 
        .C1(n7514), .Y(N28818) );
  OAI222XL U12249 ( .A0(n7475), .A1(n8002), .B0(n3515), .B1(n7999), .C0(n7513), 
        .C1(n7997), .Y(N27987) );
  OAI222XL U12250 ( .A0(n7475), .A1(n8015), .B0(n3447), .B1(n8011), .C0(n7513), 
        .C1(n8009), .Y(N28051) );
  OAI222XL U12251 ( .A0(n7475), .A1(n8027), .B0(n3378), .B1(n8024), .C0(n7513), 
        .C1(n8022), .Y(N28115) );
  OAI222XL U12252 ( .A0(n7475), .A1(n8041), .B0(n3310), .B1(n8037), .C0(n7513), 
        .C1(n8035), .Y(N28179) );
  OAI222XL U12253 ( .A0(n7475), .A1(n8079), .B0(n3097), .B1(n8075), .C0(n7513), 
        .C1(n8073), .Y(N28371) );
  OAI222XL U12254 ( .A0(n7475), .A1(n8092), .B0(n3026), .B1(n8087), .C0(n7513), 
        .C1(n8086), .Y(N28435) );
  OAI222XL U12255 ( .A0(n7475), .A1(n8155), .B0(n2543), .B1(n8152), .C0(n7513), 
        .C1(n8150), .Y(N28755) );
  OAI222XL U12256 ( .A0(n7475), .A1(n8168), .B0(n8164), .B1(n2371), .C0(n8163), 
        .C1(n7513), .Y(N28819) );
  OAI222XL U12257 ( .A0(n7477), .A1(n8015), .B0(n3446), .B1(n8012), .C0(n7512), 
        .C1(n8009), .Y(N28052) );
  OAI222XL U12258 ( .A0(n7477), .A1(n8027), .B0(n3377), .B1(n8025), .C0(n7512), 
        .C1(n8022), .Y(N28116) );
  OAI222XL U12259 ( .A0(n7477), .A1(n8079), .B0(n3096), .B1(n8075), .C0(n7512), 
        .C1(n8073), .Y(N28372) );
  OAI222XL U12260 ( .A0(n7477), .A1(n8092), .B0(n3025), .B1(n8089), .C0(n7512), 
        .C1(n8086), .Y(N28436) );
  AOI221XL U12261 ( .A0(n8509), .A1(n8158), .B0(n8510), .B1(n8147), .C0(n3915), 
        .Y(n3903) );
  OAI222XL U12262 ( .A0(n8083), .A1(n3025), .B0(n8019), .B1(n3377), .C0(n8070), 
        .C1(n3096), .Y(n3915) );
  OAI222XL U12263 ( .A0(n8518), .A1(n7933), .B0(n7930), .B1(n9000), .C0(n8004), 
        .C1(n3448), .Y(n3948) );
  OAI222XL U12264 ( .A0(n8513), .A1(n7933), .B0(n7930), .B1(n8992), .C0(n8004), 
        .C1(n3447), .Y(n3930) );
  OAI221XL U12265 ( .A0(n7473), .A1(n7990), .B0(n7514), .B1(n6591), .C0(n3586), 
        .Y(N27922) );
  OAI221XL U12266 ( .A0(n7473), .A1(n8053), .B0(n7514), .B1(n8051), .C0(n3240), 
        .Y(N28242) );
  OAI221XL U12267 ( .A0(n7473), .A1(n8103), .B0(n7514), .B1(n8102), .C0(n2957), 
        .Y(N28498) );
  OAI221XL U12268 ( .A0(n7473), .A1(n8116), .B0(n7514), .B1(n8115), .C0(n2835), 
        .Y(N28562) );
  OAI221XL U12269 ( .A0(n7473), .A1(n8130), .B0(n7514), .B1(n8128), .C0(n2750), 
        .Y(N28626) );
  OAI221XL U12270 ( .A0(n7473), .A1(n3649), .B0(n7514), .B1(n7974), .C0(n3937), 
        .Y(N27858) );
  OAI221XL U12271 ( .A0(n7475), .A1(n7990), .B0(n7513), .B1(n7987), .C0(n3585), 
        .Y(N27923) );
  OAI221XL U12272 ( .A0(n7475), .A1(n8052), .B0(n7513), .B1(n8051), .C0(n3239), 
        .Y(N28243) );
  OAI221XL U12273 ( .A0(n7475), .A1(n8103), .B0(n7513), .B1(n8102), .C0(n2956), 
        .Y(N28499) );
  OAI221XL U12274 ( .A0(n7475), .A1(n8116), .B0(n7513), .B1(n8115), .C0(n2833), 
        .Y(N28563) );
  OAI221XL U12275 ( .A0(n7475), .A1(n8130), .B0(n7513), .B1(n8128), .C0(n2749), 
        .Y(N28627) );
  OAI221XL U12276 ( .A0(n7475), .A1(n3649), .B0(n7513), .B1(n7974), .C0(n3919), 
        .Y(N27859) );
  OAI221XL U12277 ( .A0(n7477), .A1(n7990), .B0(n7512), .B1(n7987), .C0(n3584), 
        .Y(N27924) );
  AOI2BB2X1 U12278 ( .B0(n7982), .B1(n7476), .A0N(n8990), .A1N(n7979), .Y(
        n3584) );
  OAI221XL U12279 ( .A0(n7477), .A1(n8052), .B0(n7512), .B1(n8051), .C0(n3238), 
        .Y(N28244) );
  AOI2BB2X1 U12280 ( .B0(n8046), .B1(n7476), .A0N(n8988), .A1N(n8043), .Y(
        n3238) );
  OAI221XL U12281 ( .A0(n7477), .A1(n8105), .B0(n7512), .B1(n8100), .C0(n2955), 
        .Y(N28500) );
  AOI2BB2X1 U12282 ( .B0(n8098), .B1(n7476), .A0N(n8986), .A1N(n8094), .Y(
        n2955) );
  OAI221XL U12283 ( .A0(n7477), .A1(n8118), .B0(n7512), .B1(n8113), .C0(n2831), 
        .Y(N28564) );
  AOI2BB2X1 U12284 ( .B0(n8111), .B1(n7476), .A0N(n8985), .A1N(n8107), .Y(
        n2831) );
  OAI221XL U12285 ( .A0(n7477), .A1(n8131), .B0(n7512), .B1(n8126), .C0(n2748), 
        .Y(N28628) );
  AOI2BB2X1 U12286 ( .B0(n8123), .B1(n7476), .A0N(n8984), .A1N(n8120), .Y(
        n2748) );
  OAI221XL U12287 ( .A0(n7477), .A1(n3649), .B0(n7512), .B1(n7972), .C0(n3901), 
        .Y(N27860) );
  AOI2BB2X1 U12288 ( .B0(n7971), .B1(n7476), .A0N(n8983), .A1N(n7967), .Y(
        n3901) );
  OAI222XL U12289 ( .A0(n9034), .A1(n7942), .B0(n8538), .B1(n7939), .C0(n7935), 
        .C1(n9033), .Y(n4017) );
  OAI222XL U12290 ( .A0(n7958), .A1(n9031), .B0(n9038), .B1(n7955), .C0(n8538), 
        .C1(n7950), .Y(n4015) );
  OAI222XL U12291 ( .A0(n9026), .A1(n7942), .B0(n8533), .B1(n7939), .C0(n7935), 
        .C1(n9025), .Y(n3999) );
  OAI222XL U12292 ( .A0(n7956), .A1(n9023), .B0(n9030), .B1(n7955), .C0(n8533), 
        .C1(n7950), .Y(n3997) );
  OAI222XL U12293 ( .A0(n9018), .A1(n7942), .B0(n8528), .B1(n7939), .C0(n7935), 
        .C1(n9017), .Y(n3981) );
  OAI222XL U12294 ( .A0(n7957), .A1(n9015), .B0(n9022), .B1(n7955), .C0(n8528), 
        .C1(n7950), .Y(n3979) );
  OAI222XL U12295 ( .A0(n9010), .A1(n7942), .B0(n8523), .B1(n7939), .C0(n3671), 
        .C1(n9009), .Y(n3963) );
  OAI222XL U12296 ( .A0(n7958), .A1(n9007), .B0(n9014), .B1(n7955), .C0(n8523), 
        .C1(n7950), .Y(n3961) );
  OAI222XL U12297 ( .A0(n3662), .A1(n8999), .B0(n9006), .B1(n7955), .C0(n8518), 
        .C1(n7950), .Y(n3943) );
  OAI222XL U12298 ( .A0(n7463), .A1(n8002), .B0(n3521), .B1(n7999), .C0(n7519), 
        .C1(n7997), .Y(N27981) );
  OAI222XL U12299 ( .A0(n7463), .A1(n8015), .B0(n3453), .B1(n8010), .C0(n7519), 
        .C1(n8009), .Y(N28045) );
  OAI222XL U12300 ( .A0(n7463), .A1(n8028), .B0(n3384), .B1(n8024), .C0(n7519), 
        .C1(n8022), .Y(N28109) );
  OAI222XL U12301 ( .A0(n7463), .A1(n8041), .B0(n3316), .B1(n8037), .C0(n7519), 
        .C1(n8035), .Y(N28173) );
  OAI222XL U12302 ( .A0(n7463), .A1(n8079), .B0(n3103), .B1(n8075), .C0(n7519), 
        .C1(n8073), .Y(N28365) );
  OAI222XL U12303 ( .A0(n7463), .A1(n8092), .B0(n3032), .B1(n8088), .C0(n7519), 
        .C1(n8086), .Y(N28429) );
  OAI222XL U12304 ( .A0(n7463), .A1(n8155), .B0(n2549), .B1(n8152), .C0(n7519), 
        .C1(n8150), .Y(N28749) );
  OAI222XL U12305 ( .A0(n7463), .A1(n8168), .B0(n8164), .B1(n2389), .C0(n8163), 
        .C1(n7519), .Y(N28813) );
  OAI222XL U12306 ( .A0(n7465), .A1(n8002), .B0(n3520), .B1(n7999), .C0(n7518), 
        .C1(n7997), .Y(N27982) );
  OAI222XL U12307 ( .A0(n7465), .A1(n8015), .B0(n3452), .B1(n8011), .C0(n7518), 
        .C1(n8009), .Y(N28046) );
  OAI222XL U12308 ( .A0(n7465), .A1(n8028), .B0(n3383), .B1(n8024), .C0(n7518), 
        .C1(n8022), .Y(N28110) );
  OAI222XL U12309 ( .A0(n7465), .A1(n8039), .B0(n3315), .B1(n8037), .C0(n7518), 
        .C1(n8035), .Y(N28174) );
  OAI222XL U12310 ( .A0(n7465), .A1(n8079), .B0(n3102), .B1(n8075), .C0(n7518), 
        .C1(n8073), .Y(N28366) );
  OAI222XL U12311 ( .A0(n7465), .A1(n8092), .B0(n3031), .B1(n6578), .C0(n7518), 
        .C1(n8086), .Y(N28430) );
  OAI222XL U12312 ( .A0(n7465), .A1(n8155), .B0(n2548), .B1(n8152), .C0(n7518), 
        .C1(n8150), .Y(N28750) );
  OAI222XL U12313 ( .A0(n7465), .A1(n8168), .B0(n8164), .B1(n2386), .C0(n8163), 
        .C1(n7518), .Y(N28814) );
  OAI222XL U12314 ( .A0(n7467), .A1(n8002), .B0(n3519), .B1(n7999), .C0(n7517), 
        .C1(n7997), .Y(N27983) );
  OAI222XL U12315 ( .A0(n7467), .A1(n8015), .B0(n3451), .B1(n8012), .C0(n7517), 
        .C1(n8009), .Y(N28047) );
  OAI222XL U12316 ( .A0(n7467), .A1(n8028), .B0(n3382), .B1(n8025), .C0(n7517), 
        .C1(n8022), .Y(N28111) );
  OAI222XL U12317 ( .A0(n7467), .A1(n8039), .B0(n3314), .B1(n8037), .C0(n7517), 
        .C1(n8035), .Y(N28175) );
  OAI222XL U12318 ( .A0(n7467), .A1(n8079), .B0(n3101), .B1(n8075), .C0(n7517), 
        .C1(n8073), .Y(N28367) );
  OAI222XL U12319 ( .A0(n7467), .A1(n8092), .B0(n3030), .B1(n8087), .C0(n7517), 
        .C1(n8086), .Y(N28431) );
  OAI222XL U12320 ( .A0(n7467), .A1(n8155), .B0(n2547), .B1(n8152), .C0(n7517), 
        .C1(n8150), .Y(N28751) );
  OAI222XL U12321 ( .A0(n7467), .A1(n8168), .B0(n8164), .B1(n2383), .C0(n8163), 
        .C1(n7517), .Y(N28815) );
  OAI222XL U12322 ( .A0(n7469), .A1(n8002), .B0(n3518), .B1(n7999), .C0(n7516), 
        .C1(n7997), .Y(N27984) );
  OAI222XL U12323 ( .A0(n7469), .A1(n8015), .B0(n3450), .B1(n8010), .C0(n7516), 
        .C1(n8009), .Y(N28048) );
  OAI222XL U12324 ( .A0(n7469), .A1(n8028), .B0(n3381), .B1(n8023), .C0(n7516), 
        .C1(n8022), .Y(N28112) );
  OAI222XL U12325 ( .A0(n7469), .A1(n8039), .B0(n3313), .B1(n8037), .C0(n7516), 
        .C1(n8035), .Y(N28176) );
  OAI222XL U12326 ( .A0(n7469), .A1(n8079), .B0(n3100), .B1(n8075), .C0(n7516), 
        .C1(n8073), .Y(N28368) );
  OAI222XL U12327 ( .A0(n7469), .A1(n8092), .B0(n3029), .B1(n8089), .C0(n7516), 
        .C1(n8086), .Y(N28432) );
  OAI222XL U12328 ( .A0(n7469), .A1(n8155), .B0(n2546), .B1(n8152), .C0(n7516), 
        .C1(n8150), .Y(N28752) );
  OAI222XL U12329 ( .A0(n7469), .A1(n8168), .B0(n8164), .B1(n2380), .C0(n8163), 
        .C1(n7516), .Y(N28816) );
  OAI222XL U12330 ( .A0(n7471), .A1(n8002), .B0(n3517), .B1(n7999), .C0(n7515), 
        .C1(n7997), .Y(N27985) );
  OAI222XL U12331 ( .A0(n7471), .A1(n8015), .B0(n3449), .B1(n6589), .C0(n7515), 
        .C1(n8009), .Y(N28049) );
  OAI222XL U12332 ( .A0(n7471), .A1(n8028), .B0(n3380), .B1(n6577), .C0(n7515), 
        .C1(n8022), .Y(N28113) );
  OAI222XL U12333 ( .A0(n7471), .A1(n8039), .B0(n3312), .B1(n8037), .C0(n7515), 
        .C1(n8035), .Y(N28177) );
  OAI222XL U12334 ( .A0(n7471), .A1(n8079), .B0(n3099), .B1(n8075), .C0(n7515), 
        .C1(n8073), .Y(N28369) );
  OAI222XL U12335 ( .A0(n7471), .A1(n8092), .B0(n3028), .B1(n8088), .C0(n7515), 
        .C1(n8086), .Y(N28433) );
  OAI222XL U12336 ( .A0(n7471), .A1(n8155), .B0(n2545), .B1(n8152), .C0(n7515), 
        .C1(n8150), .Y(N28753) );
  OAI222XL U12337 ( .A0(n7471), .A1(n8168), .B0(n8164), .B1(n2377), .C0(n8163), 
        .C1(n7515), .Y(N28817) );
  OAI222XL U12338 ( .A0(n8543), .A1(n7933), .B0(n7930), .B1(n9040), .C0(n8004), 
        .C1(n3453), .Y(n4038) );
  OAI222XL U12339 ( .A0(n8538), .A1(n7933), .B0(n7930), .B1(n9032), .C0(n8004), 
        .C1(n3452), .Y(n4020) );
  OAI222XL U12340 ( .A0(n8533), .A1(n7933), .B0(n7930), .B1(n9024), .C0(n8006), 
        .C1(n3451), .Y(n4002) );
  OAI222XL U12341 ( .A0(n8528), .A1(n7933), .B0(n7930), .B1(n9016), .C0(n8005), 
        .C1(n3450), .Y(n3984) );
  OAI222XL U12342 ( .A0(n8523), .A1(n7933), .B0(n7930), .B1(n9008), .C0(n8006), 
        .C1(n3449), .Y(n3966) );
  OAI221XL U12343 ( .A0(n7463), .A1(n7990), .B0(n7519), .B1(n7985), .C0(n3591), 
        .Y(N27917) );
  OAI221XL U12344 ( .A0(n7463), .A1(n8052), .B0(n7519), .B1(n8050), .C0(n3245), 
        .Y(N28237) );
  OAI221XL U12345 ( .A0(n7463), .A1(n8105), .B0(n7519), .B1(n8102), .C0(n2962), 
        .Y(N28493) );
  OAI221XL U12346 ( .A0(n7463), .A1(n8118), .B0(n7519), .B1(n8115), .C0(n2845), 
        .Y(N28557) );
  OAI221XL U12347 ( .A0(n7463), .A1(n8131), .B0(n7519), .B1(n8128), .C0(n2755), 
        .Y(N28621) );
  OAI221XL U12348 ( .A0(n7463), .A1(n7977), .B0(n7519), .B1(n7974), .C0(n4027), 
        .Y(N27853) );
  OAI221XL U12349 ( .A0(n7465), .A1(n7990), .B0(n7518), .B1(n7987), .C0(n3590), 
        .Y(N27918) );
  OAI221XL U12350 ( .A0(n7465), .A1(n8052), .B0(n7518), .B1(n8049), .C0(n3244), 
        .Y(N28238) );
  OAI221XL U12351 ( .A0(n7465), .A1(n8105), .B0(n7518), .B1(n8102), .C0(n2961), 
        .Y(N28494) );
  OAI221XL U12352 ( .A0(n7465), .A1(n8118), .B0(n7518), .B1(n8115), .C0(n2843), 
        .Y(N28558) );
  OAI221XL U12353 ( .A0(n7465), .A1(n8131), .B0(n7518), .B1(n8128), .C0(n2754), 
        .Y(N28622) );
  OAI221XL U12354 ( .A0(n7465), .A1(n7976), .B0(n7518), .B1(n7974), .C0(n4009), 
        .Y(N27854) );
  OAI221XL U12355 ( .A0(n7467), .A1(n7990), .B0(n7517), .B1(n7987), .C0(n3589), 
        .Y(N27919) );
  OAI221XL U12356 ( .A0(n7467), .A1(n8052), .B0(n7517), .B1(n6592), .C0(n3243), 
        .Y(N28239) );
  OAI221XL U12357 ( .A0(n7467), .A1(n8105), .B0(n7517), .B1(n8102), .C0(n2960), 
        .Y(N28495) );
  OAI221XL U12358 ( .A0(n7467), .A1(n8118), .B0(n7517), .B1(n8115), .C0(n2841), 
        .Y(N28559) );
  OAI221XL U12359 ( .A0(n7467), .A1(n8131), .B0(n7517), .B1(n8128), .C0(n2753), 
        .Y(N28623) );
  OAI221XL U12360 ( .A0(n7467), .A1(n7977), .B0(n7517), .B1(n7974), .C0(n3991), 
        .Y(N27855) );
  OAI221XL U12361 ( .A0(n7469), .A1(n7990), .B0(n7516), .B1(n7987), .C0(n3588), 
        .Y(N27920) );
  OAI221XL U12362 ( .A0(n7469), .A1(n8052), .B0(n7516), .B1(n6592), .C0(n3242), 
        .Y(N28240) );
  OAI221XL U12363 ( .A0(n7469), .A1(n8105), .B0(n7516), .B1(n8102), .C0(n2959), 
        .Y(N28496) );
  OAI221XL U12364 ( .A0(n7469), .A1(n8118), .B0(n7516), .B1(n8115), .C0(n2839), 
        .Y(N28560) );
  OAI221XL U12365 ( .A0(n7469), .A1(n8131), .B0(n7516), .B1(n8128), .C0(n2752), 
        .Y(N28624) );
  OAI221XL U12366 ( .A0(n7469), .A1(n7977), .B0(n7516), .B1(n7974), .C0(n3973), 
        .Y(N27856) );
  OAI221XL U12367 ( .A0(n7471), .A1(n7990), .B0(n7515), .B1(n7986), .C0(n3587), 
        .Y(N27921) );
  OAI221XL U12368 ( .A0(n7471), .A1(n8053), .B0(n7515), .B1(n6592), .C0(n3241), 
        .Y(N28241) );
  OAI221XL U12369 ( .A0(n7471), .A1(n8105), .B0(n7515), .B1(n8102), .C0(n2958), 
        .Y(N28497) );
  OAI221XL U12370 ( .A0(n7471), .A1(n8118), .B0(n7515), .B1(n8115), .C0(n2837), 
        .Y(N28561) );
  OAI221XL U12371 ( .A0(n7471), .A1(n8131), .B0(n7515), .B1(n8128), .C0(n2751), 
        .Y(N28625) );
  OAI221XL U12372 ( .A0(n7471), .A1(n7977), .B0(n7515), .B1(n7974), .C0(n3955), 
        .Y(N27857) );
  OAI222XL U12373 ( .A0(n8558), .A1(n7933), .B0(n7930), .B1(n9064), .C0(n8005), 
        .C1(n3456), .Y(n4092) );
  OAI222XL U12374 ( .A0(n7958), .A1(n9063), .B0(n9070), .B1(n7954), .C0(n8558), 
        .C1(n7950), .Y(n4087) );
  OAI222XL U12375 ( .A0(n8553), .A1(n7933), .B0(n7930), .B1(n9056), .C0(n8005), 
        .C1(n3455), .Y(n4074) );
  OAI222XL U12376 ( .A0(n7957), .A1(n9055), .B0(n9062), .B1(n3663), .C0(n8553), 
        .C1(n7950), .Y(n4069) );
  OAI222XL U12377 ( .A0(n9050), .A1(n7942), .B0(n8548), .B1(n7939), .C0(n7936), 
        .C1(n9049), .Y(n4053) );
  OAI222XL U12378 ( .A0(n7957), .A1(n9047), .B0(n9054), .B1(n7954), .C0(n8548), 
        .C1(n7950), .Y(n4051) );
  OAI222XL U12379 ( .A0(n9042), .A1(n7942), .B0(n8543), .B1(n7939), .C0(n7935), 
        .C1(n9041), .Y(n4035) );
  OAI222XL U12380 ( .A0(n7957), .A1(n9039), .B0(n9046), .B1(n7954), .C0(n8543), 
        .C1(n7950), .Y(n4033) );
  OAI222XL U12381 ( .A0(n7458), .A1(n8014), .B0(n3456), .B1(n8010), .C0(n7522), 
        .C1(n8008), .Y(N28042) );
  OAI222XL U12382 ( .A0(n7458), .A1(n3362), .B0(n3387), .B1(n8023), .C0(n7522), 
        .C1(n6612), .Y(N28106) );
  OAI222XL U12383 ( .A0(n7458), .A1(n8078), .B0(n3106), .B1(n8075), .C0(n7522), 
        .C1(n8073), .Y(N28362) );
  OAI222XL U12384 ( .A0(n7458), .A1(n3010), .B0(n3035), .B1(n8087), .C0(n7522), 
        .C1(n8085), .Y(N28426) );
  OAI222XL U12385 ( .A0(n7458), .A1(n8167), .B0(n8165), .B1(n2398), .C0(n8162), 
        .C1(n7522), .Y(N28810) );
  OAI222XL U12386 ( .A0(n7460), .A1(n8014), .B0(n3455), .B1(n8011), .C0(n7521), 
        .C1(n8008), .Y(N28043) );
  OAI222XL U12387 ( .A0(n7460), .A1(n3362), .B0(n3386), .B1(n8024), .C0(n7521), 
        .C1(n8022), .Y(N28107) );
  OAI222XL U12388 ( .A0(n7460), .A1(n8078), .B0(n3105), .B1(n8075), .C0(n7521), 
        .C1(n8072), .Y(N28363) );
  OAI222XL U12389 ( .A0(n7460), .A1(n8090), .B0(n3034), .B1(n8089), .C0(n7521), 
        .C1(n8085), .Y(N28427) );
  OAI222XL U12390 ( .A0(n6623), .A1(n8015), .B0(n3454), .B1(n8012), .C0(n7520), 
        .C1(n8009), .Y(N28044) );
  OAI222XL U12391 ( .A0(n6623), .A1(n8028), .B0(n3385), .B1(n8025), .C0(n7520), 
        .C1(n8022), .Y(N28108) );
  OAI222XL U12392 ( .A0(n6623), .A1(n8079), .B0(n3104), .B1(n8075), .C0(n7520), 
        .C1(n8073), .Y(N28364) );
  OAI222XL U12393 ( .A0(n6623), .A1(n8092), .B0(n3033), .B1(n8088), .C0(n7520), 
        .C1(n8086), .Y(N28428) );
  AOI221XL U12394 ( .A0(n8559), .A1(n8159), .B0(n8560), .B1(n8146), .C0(n4095), 
        .Y(n4083) );
  OAI222XL U12395 ( .A0(n3080), .A1(n3035), .B0(n8018), .B1(n3387), .C0(n8069), 
        .C1(n3106), .Y(n4095) );
  AOI221XL U12396 ( .A0(n8554), .A1(n8159), .B0(n8555), .B1(n8146), .C0(n4077), 
        .Y(n4065) );
  OAI222XL U12397 ( .A0(n3080), .A1(n3034), .B0(n8018), .B1(n3386), .C0(n8068), 
        .C1(n3105), .Y(n4077) );
  AOI221XL U12398 ( .A0(n8549), .A1(n8159), .B0(n8550), .B1(n8147), .C0(n4059), 
        .Y(n4047) );
  OAI222XL U12399 ( .A0(n8080), .A1(n3033), .B0(n8018), .B1(n3385), .C0(n8068), 
        .C1(n3104), .Y(n4059) );
  AOI221XL U12400 ( .A0(n8551), .A1(n7991), .B0(n8552), .B1(n8032), .C0(n4056), 
        .Y(n4048) );
  OAI222XL U12401 ( .A0(n8548), .A1(n7933), .B0(n7930), .B1(n9048), .C0(n8004), 
        .C1(n3454), .Y(n4056) );
  OAI221XL U12402 ( .A0(n7458), .A1(n7990), .B0(n7522), .B1(n6591), .C0(n3594), 
        .Y(N27914) );
  OAI221XL U12403 ( .A0(n7458), .A1(n8053), .B0(n7522), .B1(n6592), .C0(n3248), 
        .Y(N28234) );
  AOI2BB2X1 U12404 ( .B0(n8047), .B1(n7457), .A0N(n9068), .A1N(n8043), .Y(
        n3248) );
  OAI221XL U12405 ( .A0(n7458), .A1(n8103), .B0(n7522), .B1(n8102), .C0(n2965), 
        .Y(N28490) );
  OAI221XL U12406 ( .A0(n7458), .A1(n8116), .B0(n7522), .B1(n8115), .C0(n2851), 
        .Y(N28554) );
  OAI221XL U12407 ( .A0(n7458), .A1(n8130), .B0(n7522), .B1(n8128), .C0(n2758), 
        .Y(N28618) );
  OAI221XL U12408 ( .A0(n7458), .A1(n3649), .B0(n7522), .B1(n7974), .C0(n4081), 
        .Y(N27850) );
  OAI221XL U12409 ( .A0(n7460), .A1(n7990), .B0(n7521), .B1(n7985), .C0(n3593), 
        .Y(N27915) );
  AOI2BB2X1 U12410 ( .B0(n7983), .B1(n7459), .A0N(n9062), .A1N(n7979), .Y(
        n3593) );
  OAI221XL U12411 ( .A0(n7460), .A1(n8053), .B0(n7521), .B1(n6592), .C0(n3247), 
        .Y(N28235) );
  AOI2BB2X1 U12412 ( .B0(n8047), .B1(n7459), .A0N(n9060), .A1N(n8043), .Y(
        n3247) );
  OAI221XL U12413 ( .A0(n7460), .A1(n8105), .B0(n7521), .B1(n8102), .C0(n2964), 
        .Y(N28491) );
  AOI2BB2X1 U12414 ( .B0(n8099), .B1(n7459), .A0N(n9058), .A1N(n8094), .Y(
        n2964) );
  OAI221XL U12415 ( .A0(n7460), .A1(n8116), .B0(n7521), .B1(n8115), .C0(n2849), 
        .Y(N28555) );
  AOI2BB2X1 U12416 ( .B0(n8112), .B1(n7459), .A0N(n9057), .A1N(n8107), .Y(
        n2849) );
  OAI221XL U12417 ( .A0(n7460), .A1(n8131), .B0(n7521), .B1(n8128), .C0(n2757), 
        .Y(N28619) );
  AOI2BB2X1 U12418 ( .B0(n8124), .B1(n7459), .A0N(n9056), .A1N(n8120), .Y(
        n2757) );
  OAI221XL U12419 ( .A0(n7460), .A1(n7977), .B0(n7521), .B1(n7974), .C0(n4063), 
        .Y(N27851) );
  AOI2BB2X1 U12420 ( .B0(n7969), .B1(n7459), .A0N(n9055), .A1N(n7967), .Y(
        n4063) );
  OAI221XL U12421 ( .A0(n6623), .A1(n7990), .B0(n7520), .B1(n6591), .C0(n3592), 
        .Y(N27916) );
  AOI2BB2X1 U12422 ( .B0(n7983), .B1(n7461), .A0N(n9054), .A1N(n7979), .Y(
        n3592) );
  OAI221XL U12423 ( .A0(n6623), .A1(n8053), .B0(n7520), .B1(n6592), .C0(n3246), 
        .Y(N28236) );
  AOI2BB2X1 U12424 ( .B0(n8047), .B1(n7461), .A0N(n9052), .A1N(n8043), .Y(
        n3246) );
  OAI221XL U12425 ( .A0(n6623), .A1(n8103), .B0(n7520), .B1(n8102), .C0(n2963), 
        .Y(N28492) );
  AOI2BB2X1 U12426 ( .B0(n8099), .B1(n7461), .A0N(n9050), .A1N(n8094), .Y(
        n2963) );
  OAI221XL U12427 ( .A0(n6623), .A1(n8116), .B0(n7520), .B1(n8115), .C0(n2847), 
        .Y(N28556) );
  AOI2BB2X1 U12428 ( .B0(n8112), .B1(n7461), .A0N(n9049), .A1N(n8107), .Y(
        n2847) );
  OAI221XL U12429 ( .A0(n6623), .A1(n8131), .B0(n7520), .B1(n8128), .C0(n2756), 
        .Y(N28620) );
  AOI2BB2X1 U12430 ( .B0(n8125), .B1(n7461), .A0N(n9048), .A1N(n8120), .Y(
        n2756) );
  OAI221XL U12431 ( .A0(n6623), .A1(n7977), .B0(n7520), .B1(n7974), .C0(n4045), 
        .Y(N27852) );
  AOI2BB2X1 U12432 ( .B0(n7969), .B1(n7461), .A0N(n9047), .A1N(n7967), .Y(
        n4045) );
  OAI222XL U12433 ( .A0(n9098), .A1(n3669), .B0(n8578), .B1(n7940), .C0(n7937), 
        .C1(n9097), .Y(n4161) );
  OAI222XL U12434 ( .A0(n7957), .A1(n9095), .B0(n9102), .B1(n7953), .C0(n8578), 
        .C1(n7951), .Y(n4159) );
  OAI222XL U12435 ( .A0(n9090), .A1(n7943), .B0(n8573), .B1(n7940), .C0(n7936), 
        .C1(n9089), .Y(n4143) );
  OAI222XL U12436 ( .A0(n7958), .A1(n9087), .B0(n9094), .B1(n7953), .C0(n8573), 
        .C1(n7951), .Y(n4141) );
  OAI222XL U12437 ( .A0(n9082), .A1(n7941), .B0(n8568), .B1(n7940), .C0(n7935), 
        .C1(n9081), .Y(n4125) );
  OAI222XL U12438 ( .A0(n3662), .A1(n9079), .B0(n9086), .B1(n7953), .C0(n8568), 
        .C1(n7951), .Y(n4123) );
  OAI222XL U12439 ( .A0(n9074), .A1(n7942), .B0(n8563), .B1(n7939), .C0(n7936), 
        .C1(n9073), .Y(n4107) );
  OAI222XL U12440 ( .A0(n3662), .A1(n9071), .B0(n9078), .B1(n7955), .C0(n8563), 
        .C1(n7950), .Y(n4105) );
  OAI222XL U12441 ( .A0(n7448), .A1(n8003), .B0(n3529), .B1(n8000), .C0(n7527), 
        .C1(n7996), .Y(N27973) );
  OAI222XL U12442 ( .A0(n7448), .A1(n8014), .B0(n3461), .B1(n8011), .C0(n7527), 
        .C1(n8008), .Y(N28037) );
  OAI222XL U12443 ( .A0(n7448), .A1(n8028), .B0(n3392), .B1(n8024), .C0(n7527), 
        .C1(n8021), .Y(N28101) );
  OAI222XL U12444 ( .A0(n7448), .A1(n8041), .B0(n3324), .B1(n8038), .C0(n7527), 
        .C1(n8035), .Y(N28165) );
  OAI222XL U12445 ( .A0(n7448), .A1(n8078), .B0(n3111), .B1(n8076), .C0(n7527), 
        .C1(n8073), .Y(N28357) );
  OAI222XL U12446 ( .A0(n7448), .A1(n8092), .B0(n3040), .B1(n8088), .C0(n7527), 
        .C1(n8085), .Y(N28421) );
  OAI222XL U12447 ( .A0(n7448), .A1(n8156), .B0(n2557), .B1(n8153), .C0(n7527), 
        .C1(n8149), .Y(N28741) );
  OAI222XL U12448 ( .A0(n7448), .A1(n8167), .B0(n8166), .B1(n2413), .C0(n8161), 
        .C1(n7527), .Y(N28805) );
  OAI222XL U12449 ( .A0(n7450), .A1(n8003), .B0(n3528), .B1(n8000), .C0(n7526), 
        .C1(n7996), .Y(N27974) );
  OAI222XL U12450 ( .A0(n7450), .A1(n8014), .B0(n3460), .B1(n8011), .C0(n7526), 
        .C1(n8008), .Y(N28038) );
  OAI222XL U12451 ( .A0(n7450), .A1(n8027), .B0(n3391), .B1(n8024), .C0(n7526), 
        .C1(n8022), .Y(N28102) );
  OAI222XL U12452 ( .A0(n7450), .A1(n8040), .B0(n3323), .B1(n8038), .C0(n7526), 
        .C1(n8033), .Y(N28166) );
  OAI222XL U12453 ( .A0(n7450), .A1(n8078), .B0(n3110), .B1(n8076), .C0(n7526), 
        .C1(n8073), .Y(N28358) );
  OAI222XL U12454 ( .A0(n7450), .A1(n8091), .B0(n3039), .B1(n8088), .C0(n7526), 
        .C1(n8085), .Y(N28422) );
  OAI222XL U12455 ( .A0(n7450), .A1(n8156), .B0(n2556), .B1(n8153), .C0(n7526), 
        .C1(n8149), .Y(N28742) );
  OAI222XL U12456 ( .A0(n7450), .A1(n8167), .B0(n8166), .B1(n2410), .C0(n6616), 
        .C1(n7526), .Y(N28806) );
  OAI222XL U12457 ( .A0(n7452), .A1(n8003), .B0(n3527), .B1(n8000), .C0(n7525), 
        .C1(n7996), .Y(N27975) );
  OAI222XL U12458 ( .A0(n7452), .A1(n8014), .B0(n3459), .B1(n8011), .C0(n7525), 
        .C1(n8008), .Y(N28039) );
  OAI222XL U12459 ( .A0(n7452), .A1(n8028), .B0(n3390), .B1(n8024), .C0(n7525), 
        .C1(n8022), .Y(N28103) );
  OAI222XL U12460 ( .A0(n7452), .A1(n8040), .B0(n3322), .B1(n8038), .C0(n7525), 
        .C1(n8033), .Y(N28167) );
  OAI222XL U12461 ( .A0(n7452), .A1(n8078), .B0(n3109), .B1(n8076), .C0(n7525), 
        .C1(n8073), .Y(N28359) );
  OAI222XL U12462 ( .A0(n7452), .A1(n8092), .B0(n3038), .B1(n8088), .C0(n7525), 
        .C1(n8085), .Y(N28423) );
  OAI222XL U12463 ( .A0(n7452), .A1(n8156), .B0(n2555), .B1(n8153), .C0(n7525), 
        .C1(n8149), .Y(N28743) );
  OAI222XL U12464 ( .A0(n7452), .A1(n8167), .B0(n8164), .B1(n2407), .C0(n8163), 
        .C1(n7525), .Y(N28807) );
  OAI222XL U12465 ( .A0(n7454), .A1(n8003), .B0(n3526), .B1(n8000), .C0(n7524), 
        .C1(n7996), .Y(N27976) );
  OAI222XL U12466 ( .A0(n7454), .A1(n8014), .B0(n3458), .B1(n8011), .C0(n7524), 
        .C1(n8008), .Y(N28040) );
  OAI222XL U12467 ( .A0(n7454), .A1(n8028), .B0(n3389), .B1(n8024), .C0(n7524), 
        .C1(n8022), .Y(N28104) );
  OAI222XL U12468 ( .A0(n7454), .A1(n8040), .B0(n3321), .B1(n8038), .C0(n7524), 
        .C1(n6613), .Y(N28168) );
  OAI222XL U12469 ( .A0(n7454), .A1(n8078), .B0(n3108), .B1(n8076), .C0(n7524), 
        .C1(n8073), .Y(N28360) );
  OAI222XL U12470 ( .A0(n7454), .A1(n8092), .B0(n3037), .B1(n8088), .C0(n7524), 
        .C1(n8085), .Y(N28424) );
  OAI222XL U12471 ( .A0(n7454), .A1(n8156), .B0(n2554), .B1(n8153), .C0(n7524), 
        .C1(n8149), .Y(N28744) );
  OAI222XL U12472 ( .A0(n7454), .A1(n8167), .B0(n8165), .B1(n2404), .C0(n6616), 
        .C1(n7524), .Y(N28808) );
  OAI222XL U12473 ( .A0(n7456), .A1(n8001), .B0(n3525), .B1(n7999), .C0(n7523), 
        .C1(n7996), .Y(N27977) );
  OAI222XL U12474 ( .A0(n7456), .A1(n8014), .B0(n3457), .B1(n8012), .C0(n7523), 
        .C1(n8008), .Y(N28041) );
  OAI222XL U12475 ( .A0(n7456), .A1(n8026), .B0(n3388), .B1(n8025), .C0(n7523), 
        .C1(n8020), .Y(N28105) );
  OAI222XL U12476 ( .A0(n7456), .A1(n8041), .B0(n3320), .B1(n8037), .C0(n7523), 
        .C1(n6613), .Y(N28169) );
  OAI222XL U12477 ( .A0(n7456), .A1(n8078), .B0(n3107), .B1(n8075), .C0(n7523), 
        .C1(n8071), .Y(N28361) );
  OAI222XL U12478 ( .A0(n7456), .A1(n8090), .B0(n3036), .B1(n8087), .C0(n7523), 
        .C1(n8085), .Y(N28425) );
  OAI222XL U12479 ( .A0(n7456), .A1(n8156), .B0(n2553), .B1(n8152), .C0(n7523), 
        .C1(n8149), .Y(N28745) );
  OAI222XL U12480 ( .A0(n7456), .A1(n8167), .B0(n8165), .B1(n2401), .C0(n6616), 
        .C1(n7523), .Y(N28809) );
  OAI222XL U12481 ( .A0(n8583), .A1(n7934), .B0(n7931), .B1(n9104), .C0(n8006), 
        .C1(n3461), .Y(n4182) );
  OAI222XL U12482 ( .A0(n8578), .A1(n7934), .B0(n7931), .B1(n9096), .C0(n8006), 
        .C1(n3460), .Y(n4164) );
  OAI222XL U12483 ( .A0(n8573), .A1(n7934), .B0(n7930), .B1(n9088), .C0(n8004), 
        .C1(n3459), .Y(n4146) );
  OAI222XL U12484 ( .A0(n8568), .A1(n7934), .B0(n7930), .B1(n9080), .C0(n8004), 
        .C1(n3458), .Y(n4128) );
  OAI222XL U12485 ( .A0(n8563), .A1(n7933), .B0(n7930), .B1(n9072), .C0(n8004), 
        .C1(n3457), .Y(n4110) );
  OAI221XL U12486 ( .A0(n7448), .A1(n7988), .B0(n7527), .B1(n6591), .C0(n3599), 
        .Y(N27909) );
  OAI221XL U12487 ( .A0(n7448), .A1(n8054), .B0(n7527), .B1(n8049), .C0(n3253), 
        .Y(N28229) );
  OAI221XL U12488 ( .A0(n7448), .A1(n8103), .B0(n7527), .B1(n6599), .C0(n2970), 
        .Y(N28485) );
  OAI221XL U12489 ( .A0(n7448), .A1(n8118), .B0(n7527), .B1(n6598), .C0(n2861), 
        .Y(N28549) );
  OAI221XL U12490 ( .A0(n7448), .A1(n6609), .B0(n7527), .B1(n6600), .C0(n2763), 
        .Y(N28613) );
  OAI221XL U12491 ( .A0(n7448), .A1(n7977), .B0(n7527), .B1(n7973), .C0(n4171), 
        .Y(N27845) );
  OAI221XL U12492 ( .A0(n7450), .A1(n7989), .B0(n7526), .B1(n7987), .C0(n3598), 
        .Y(N27910) );
  OAI221XL U12493 ( .A0(n7450), .A1(n8054), .B0(n7526), .B1(n8049), .C0(n3252), 
        .Y(N28230) );
  OAI221XL U12494 ( .A0(n7450), .A1(n8103), .B0(n7526), .B1(n6599), .C0(n2969), 
        .Y(N28486) );
  OAI221XL U12495 ( .A0(n7450), .A1(n8118), .B0(n7526), .B1(n6598), .C0(n2859), 
        .Y(N28550) );
  OAI221XL U12496 ( .A0(n7450), .A1(n8129), .B0(n7526), .B1(n8126), .C0(n2762), 
        .Y(N28614) );
  OAI221XL U12497 ( .A0(n7450), .A1(n7977), .B0(n7526), .B1(n7974), .C0(n4153), 
        .Y(N27846) );
  OAI221XL U12498 ( .A0(n7452), .A1(n7989), .B0(n7525), .B1(n7985), .C0(n3597), 
        .Y(N27911) );
  OAI221XL U12499 ( .A0(n7452), .A1(n8054), .B0(n7525), .B1(n8049), .C0(n3251), 
        .Y(N28231) );
  OAI221XL U12500 ( .A0(n7452), .A1(n8104), .B0(n7525), .B1(n8102), .C0(n2968), 
        .Y(N28487) );
  OAI221XL U12501 ( .A0(n7452), .A1(n8118), .B0(n7525), .B1(n8115), .C0(n2857), 
        .Y(N28551) );
  OAI221XL U12502 ( .A0(n7452), .A1(n8129), .B0(n7525), .B1(n8128), .C0(n2761), 
        .Y(N28615) );
  OAI221XL U12503 ( .A0(n7452), .A1(n7977), .B0(n7525), .B1(n7974), .C0(n4135), 
        .Y(N27847) );
  OAI221XL U12504 ( .A0(n7454), .A1(n7989), .B0(n7524), .B1(n7985), .C0(n3596), 
        .Y(N27912) );
  OAI221XL U12505 ( .A0(n7454), .A1(n8054), .B0(n7524), .B1(n8049), .C0(n3250), 
        .Y(N28232) );
  OAI221XL U12506 ( .A0(n7454), .A1(n8104), .B0(n7524), .B1(n8102), .C0(n2967), 
        .Y(N28488) );
  OAI221XL U12507 ( .A0(n7454), .A1(n8118), .B0(n7524), .B1(n8115), .C0(n2855), 
        .Y(N28552) );
  OAI221XL U12508 ( .A0(n7454), .A1(n8129), .B0(n7524), .B1(n8128), .C0(n2760), 
        .Y(N28616) );
  OAI221XL U12509 ( .A0(n7454), .A1(n7977), .B0(n7524), .B1(n7974), .C0(n4117), 
        .Y(N27848) );
  OAI221XL U12510 ( .A0(n7456), .A1(n7990), .B0(n7523), .B1(n7985), .C0(n3595), 
        .Y(N27913) );
  OAI221XL U12511 ( .A0(n7456), .A1(n8053), .B0(n7523), .B1(n8049), .C0(n3249), 
        .Y(N28233) );
  OAI221XL U12512 ( .A0(n7456), .A1(n8105), .B0(n7523), .B1(n8102), .C0(n2966), 
        .Y(N28489) );
  OAI221XL U12513 ( .A0(n7456), .A1(n8118), .B0(n7523), .B1(n8115), .C0(n2853), 
        .Y(N28553) );
  OAI221XL U12514 ( .A0(n7456), .A1(n8130), .B0(n7523), .B1(n8128), .C0(n2759), 
        .Y(N28617) );
  OAI221XL U12515 ( .A0(n7456), .A1(n3649), .B0(n7523), .B1(n7974), .C0(n4099), 
        .Y(N27849) );
  OAI222XL U12516 ( .A0(n8603), .A1(n7934), .B0(n7931), .B1(n9136), .C0(n8005), 
        .C1(n3465), .Y(n4254) );
  OAI222XL U12517 ( .A0(n7957), .A1(n9135), .B0(n9142), .B1(n7953), .C0(n8603), 
        .C1(n7951), .Y(n4249) );
  OAI222XL U12518 ( .A0(n9130), .A1(n7942), .B0(n8598), .B1(n7940), .C0(n7937), 
        .C1(n9129), .Y(n4233) );
  OAI222XL U12519 ( .A0(n7957), .A1(n9127), .B0(n9134), .B1(n7953), .C0(n8598), 
        .C1(n7951), .Y(n4231) );
  OAI222XL U12520 ( .A0(n9122), .A1(n7941), .B0(n8593), .B1(n7940), .C0(n7937), 
        .C1(n9121), .Y(n4215) );
  OAI222XL U12521 ( .A0(n7957), .A1(n9119), .B0(n9126), .B1(n7953), .C0(n8593), 
        .C1(n7951), .Y(n4213) );
  OAI222XL U12522 ( .A0(n9114), .A1(n7942), .B0(n8588), .B1(n7940), .C0(n7937), 
        .C1(n9113), .Y(n4197) );
  OAI222XL U12523 ( .A0(n7957), .A1(n9111), .B0(n9118), .B1(n7953), .C0(n8588), 
        .C1(n7951), .Y(n4195) );
  OAI222XL U12524 ( .A0(n9106), .A1(n3669), .B0(n8583), .B1(n7940), .C0(n7937), 
        .C1(n9105), .Y(n4179) );
  OAI222XL U12525 ( .A0(n7957), .A1(n9103), .B0(n9110), .B1(n7953), .C0(n8583), 
        .C1(n7951), .Y(n4177) );
  OAI222XL U12526 ( .A0(n7440), .A1(n8014), .B0(n3465), .B1(n8011), .C0(n7531), 
        .C1(n8008), .Y(N28033) );
  OAI222XL U12527 ( .A0(n7440), .A1(n8026), .B0(n3396), .B1(n8024), .C0(n7531), 
        .C1(n8020), .Y(N28097) );
  OAI222XL U12528 ( .A0(n7440), .A1(n8078), .B0(n3115), .B1(n8076), .C0(n7531), 
        .C1(n8071), .Y(N28353) );
  OAI222XL U12529 ( .A0(n7440), .A1(n8092), .B0(n3044), .B1(n8088), .C0(n7531), 
        .C1(n8085), .Y(N28417) );
  OAI222XL U12530 ( .A0(n7440), .A1(n8167), .B0(n8166), .B1(n2425), .C0(n6616), 
        .C1(n7531), .Y(N28801) );
  OAI222XL U12531 ( .A0(n7442), .A1(n8003), .B0(n3532), .B1(n8000), .C0(n7530), 
        .C1(n7996), .Y(N27970) );
  OAI222XL U12532 ( .A0(n7442), .A1(n8014), .B0(n3464), .B1(n8011), .C0(n7530), 
        .C1(n8008), .Y(N28034) );
  OAI222XL U12533 ( .A0(n7442), .A1(n8028), .B0(n3395), .B1(n8024), .C0(n7530), 
        .C1(n8022), .Y(N28098) );
  OAI222XL U12534 ( .A0(n7442), .A1(n8040), .B0(n3327), .B1(n8038), .C0(n7530), 
        .C1(n6613), .Y(N28162) );
  OAI222XL U12535 ( .A0(n7442), .A1(n8078), .B0(n3114), .B1(n8076), .C0(n7530), 
        .C1(n8071), .Y(N28354) );
  OAI222XL U12536 ( .A0(n7442), .A1(n8092), .B0(n3043), .B1(n8088), .C0(n7530), 
        .C1(n8085), .Y(N28418) );
  OAI222XL U12537 ( .A0(n7442), .A1(n8156), .B0(n2560), .B1(n8153), .C0(n7530), 
        .C1(n8149), .Y(N28738) );
  OAI222XL U12538 ( .A0(n7442), .A1(n8167), .B0(n8166), .B1(n2422), .C0(n6616), 
        .C1(n7530), .Y(N28802) );
  OAI222XL U12539 ( .A0(n7444), .A1(n8003), .B0(n3531), .B1(n8000), .C0(n7529), 
        .C1(n7996), .Y(N27971) );
  OAI222XL U12540 ( .A0(n7444), .A1(n8014), .B0(n3463), .B1(n8011), .C0(n7529), 
        .C1(n8008), .Y(N28035) );
  OAI222XL U12541 ( .A0(n7444), .A1(n8028), .B0(n3394), .B1(n8024), .C0(n7529), 
        .C1(n8020), .Y(N28099) );
  OAI222XL U12542 ( .A0(n7444), .A1(n8040), .B0(n3326), .B1(n8038), .C0(n7529), 
        .C1(n6613), .Y(N28163) );
  OAI222XL U12543 ( .A0(n7444), .A1(n8078), .B0(n3113), .B1(n8076), .C0(n7529), 
        .C1(n6614), .Y(N28355) );
  OAI222XL U12544 ( .A0(n7444), .A1(n8090), .B0(n3042), .B1(n8088), .C0(n7529), 
        .C1(n8085), .Y(N28419) );
  OAI222XL U12545 ( .A0(n7444), .A1(n8154), .B0(n2559), .B1(n8153), .C0(n7529), 
        .C1(n8149), .Y(N28739) );
  OAI222XL U12546 ( .A0(n7444), .A1(n8167), .B0(n8166), .B1(n2419), .C0(n6616), 
        .C1(n7529), .Y(N28803) );
  OAI222XL U12547 ( .A0(n7446), .A1(n8003), .B0(n3530), .B1(n8000), .C0(n7528), 
        .C1(n7996), .Y(N27972) );
  OAI222XL U12548 ( .A0(n7446), .A1(n8014), .B0(n3462), .B1(n8011), .C0(n7528), 
        .C1(n8008), .Y(N28036) );
  OAI222XL U12549 ( .A0(n7446), .A1(n8026), .B0(n3393), .B1(n8024), .C0(n7528), 
        .C1(n8020), .Y(N28100) );
  OAI222XL U12550 ( .A0(n7446), .A1(n8040), .B0(n3325), .B1(n8038), .C0(n7528), 
        .C1(n6613), .Y(N28164) );
  OAI222XL U12551 ( .A0(n7446), .A1(n8078), .B0(n3112), .B1(n8076), .C0(n7528), 
        .C1(n6614), .Y(N28356) );
  OAI222XL U12552 ( .A0(n7446), .A1(n8090), .B0(n3041), .B1(n8088), .C0(n7528), 
        .C1(n8085), .Y(N28420) );
  OAI222XL U12553 ( .A0(n7446), .A1(n8154), .B0(n2558), .B1(n8153), .C0(n7528), 
        .C1(n8149), .Y(N28740) );
  OAI222XL U12554 ( .A0(n7446), .A1(n8167), .B0(n8166), .B1(n2416), .C0(n8163), 
        .C1(n7528), .Y(N28804) );
  AOI221XL U12555 ( .A0(n8604), .A1(n8160), .B0(n8605), .B1(n8146), .C0(n4257), 
        .Y(n4245) );
  OAI222XL U12556 ( .A0(n8082), .A1(n3044), .B0(n8018), .B1(n3396), .C0(n8069), 
        .C1(n3115), .Y(n4257) );
  OAI222XL U12557 ( .A0(n8598), .A1(n7934), .B0(n7931), .B1(n9128), .C0(n8006), 
        .C1(n3464), .Y(n4236) );
  OAI222XL U12558 ( .A0(n8593), .A1(n7934), .B0(n7931), .B1(n9120), .C0(n3498), 
        .C1(n3463), .Y(n4218) );
  OAI222XL U12559 ( .A0(n8588), .A1(n7934), .B0(n7931), .B1(n9112), .C0(n3498), 
        .C1(n3462), .Y(n4200) );
  OAI221XL U12560 ( .A0(n7440), .A1(n7988), .B0(n7531), .B1(n6591), .C0(n3603), 
        .Y(N27905) );
  OAI221XL U12561 ( .A0(n7440), .A1(n8054), .B0(n7531), .B1(n8049), .C0(n3257), 
        .Y(N28225) );
  AOI2BB2X1 U12562 ( .B0(n8048), .B1(n7439), .A0N(n9140), .A1N(n8044), .Y(
        n3257) );
  OAI221XL U12563 ( .A0(n7440), .A1(n8105), .B0(n7531), .B1(n8100), .C0(n2974), 
        .Y(N28481) );
  OAI221XL U12564 ( .A0(n7440), .A1(n8118), .B0(n7531), .B1(n6598), .C0(n2869), 
        .Y(N28545) );
  OAI221XL U12565 ( .A0(n7440), .A1(n8130), .B0(n7531), .B1(n8126), .C0(n2767), 
        .Y(N28609) );
  OAI221XL U12566 ( .A0(n7440), .A1(n7977), .B0(n7531), .B1(n7973), .C0(n4243), 
        .Y(N27841) );
  OAI221XL U12567 ( .A0(n7442), .A1(n7989), .B0(n7530), .B1(n7987), .C0(n3602), 
        .Y(N27906) );
  OAI221XL U12568 ( .A0(n7442), .A1(n8054), .B0(n7530), .B1(n8049), .C0(n3256), 
        .Y(N28226) );
  OAI221XL U12569 ( .A0(n7442), .A1(n8103), .B0(n7530), .B1(n6599), .C0(n2973), 
        .Y(N28482) );
  OAI221XL U12570 ( .A0(n7442), .A1(n8118), .B0(n7530), .B1(n8115), .C0(n2867), 
        .Y(N28546) );
  OAI221XL U12571 ( .A0(n7442), .A1(n8131), .B0(n7530), .B1(n8128), .C0(n2766), 
        .Y(N28610) );
  OAI221XL U12572 ( .A0(n7442), .A1(n7977), .B0(n7530), .B1(n7974), .C0(n4225), 
        .Y(N27842) );
  OAI221XL U12573 ( .A0(n7444), .A1(n7988), .B0(n7529), .B1(n6591), .C0(n3601), 
        .Y(N27907) );
  OAI221XL U12574 ( .A0(n7444), .A1(n8054), .B0(n7529), .B1(n8050), .C0(n3255), 
        .Y(N28227) );
  OAI221XL U12575 ( .A0(n7444), .A1(n8104), .B0(n7529), .B1(n8100), .C0(n2972), 
        .Y(N28483) );
  OAI221XL U12576 ( .A0(n7444), .A1(n8118), .B0(n7529), .B1(n8113), .C0(n2865), 
        .Y(N28547) );
  OAI221XL U12577 ( .A0(n7444), .A1(n6609), .B0(n7529), .B1(n6600), .C0(n2765), 
        .Y(N28611) );
  OAI221XL U12578 ( .A0(n7444), .A1(n7977), .B0(n7529), .B1(n7974), .C0(n4207), 
        .Y(N27843) );
  OAI221XL U12579 ( .A0(n7446), .A1(n7989), .B0(n7528), .B1(n7987), .C0(n3600), 
        .Y(N27908) );
  OAI221XL U12580 ( .A0(n7446), .A1(n8054), .B0(n7528), .B1(n8051), .C0(n3254), 
        .Y(N28228) );
  OAI221XL U12581 ( .A0(n7446), .A1(n8104), .B0(n7528), .B1(n8100), .C0(n2971), 
        .Y(N28484) );
  OAI221XL U12582 ( .A0(n7446), .A1(n8118), .B0(n7528), .B1(n8113), .C0(n2863), 
        .Y(N28548) );
  OAI221XL U12583 ( .A0(n7446), .A1(n8129), .B0(n7528), .B1(n8126), .C0(n2764), 
        .Y(N28612) );
  OAI221XL U12584 ( .A0(n7446), .A1(n7977), .B0(n7528), .B1(n7974), .C0(n4189), 
        .Y(N27844) );
  OAI222XL U12585 ( .A0(n9162), .A1(n7941), .B0(n8618), .B1(n7940), .C0(n7937), 
        .C1(n9161), .Y(n4305) );
  OAI222XL U12586 ( .A0(n7957), .A1(n9159), .B0(n9166), .B1(n7953), .C0(n8618), 
        .C1(n7951), .Y(n4303) );
  OAI222XL U12587 ( .A0(n9154), .A1(n7942), .B0(n8613), .B1(n7940), .C0(n7937), 
        .C1(n9153), .Y(n4287) );
  OAI222XL U12588 ( .A0(n7957), .A1(n9151), .B0(n9158), .B1(n7953), .C0(n8613), 
        .C1(n7951), .Y(n4285) );
  OAI222XL U12589 ( .A0(n8608), .A1(n7934), .B0(n7931), .B1(n9144), .C0(n8005), 
        .C1(n3466), .Y(n4272) );
  OAI222XL U12590 ( .A0(n7957), .A1(n9143), .B0(n9150), .B1(n7953), .C0(n8608), 
        .C1(n7951), .Y(n4267) );
  OAI222XL U12591 ( .A0(n7432), .A1(n8003), .B0(n3537), .B1(n8000), .C0(n7535), 
        .C1(n7996), .Y(N27965) );
  OAI222XL U12592 ( .A0(n7432), .A1(n8014), .B0(n3469), .B1(n8011), .C0(n7535), 
        .C1(n8008), .Y(N28029) );
  OAI222XL U12593 ( .A0(n7432), .A1(n8026), .B0(n3400), .B1(n8024), .C0(n7535), 
        .C1(n6612), .Y(N28093) );
  OAI222XL U12594 ( .A0(n7432), .A1(n8041), .B0(n3332), .B1(n8038), .C0(n7535), 
        .C1(n6613), .Y(N28157) );
  OAI222XL U12595 ( .A0(n7432), .A1(n8078), .B0(n3119), .B1(n8076), .C0(n7535), 
        .C1(n6614), .Y(N28349) );
  OAI222XL U12596 ( .A0(n7432), .A1(n8090), .B0(n3048), .B1(n8088), .C0(n7535), 
        .C1(n8085), .Y(N28413) );
  OAI222XL U12597 ( .A0(n7432), .A1(n8154), .B0(n2565), .B1(n8153), .C0(n7535), 
        .C1(n8149), .Y(N28733) );
  OAI222XL U12598 ( .A0(n7432), .A1(n8167), .B0(n8166), .B1(n2437), .C0(n8161), 
        .C1(n7535), .Y(N28797) );
  OAI222XL U12599 ( .A0(n7434), .A1(n8003), .B0(n3536), .B1(n8000), .C0(n7534), 
        .C1(n7996), .Y(N27966) );
  OAI222XL U12600 ( .A0(n7434), .A1(n8014), .B0(n3468), .B1(n8011), .C0(n7534), 
        .C1(n8008), .Y(N28030) );
  OAI222XL U12601 ( .A0(n7434), .A1(n8026), .B0(n3399), .B1(n8024), .C0(n7534), 
        .C1(n6612), .Y(N28094) );
  OAI222XL U12602 ( .A0(n7434), .A1(n8041), .B0(n3331), .B1(n8038), .C0(n7534), 
        .C1(n8033), .Y(N28158) );
  OAI222XL U12603 ( .A0(n7434), .A1(n8078), .B0(n3118), .B1(n8076), .C0(n7534), 
        .C1(n6614), .Y(N28350) );
  OAI222XL U12604 ( .A0(n7434), .A1(n3010), .B0(n3047), .B1(n8088), .C0(n7534), 
        .C1(n8085), .Y(N28414) );
  OAI222XL U12605 ( .A0(n7434), .A1(n8154), .B0(n2564), .B1(n8153), .C0(n7534), 
        .C1(n8149), .Y(N28734) );
  OAI222XL U12606 ( .A0(n7434), .A1(n8167), .B0(n8166), .B1(n2434), .C0(n8163), 
        .C1(n7534), .Y(N28798) );
  OAI222XL U12607 ( .A0(n7436), .A1(n8003), .B0(n3535), .B1(n8000), .C0(n7533), 
        .C1(n7996), .Y(N27967) );
  OAI222XL U12608 ( .A0(n7436), .A1(n8014), .B0(n3467), .B1(n8011), .C0(n7533), 
        .C1(n8008), .Y(N28031) );
  OAI222XL U12609 ( .A0(n7436), .A1(n3362), .B0(n3398), .B1(n8024), .C0(n7533), 
        .C1(n6612), .Y(N28095) );
  OAI222XL U12610 ( .A0(n7436), .A1(n6576), .B0(n3330), .B1(n8038), .C0(n7533), 
        .C1(n8033), .Y(N28159) );
  OAI222XL U12611 ( .A0(n7436), .A1(n8078), .B0(n3117), .B1(n8076), .C0(n7533), 
        .C1(n6614), .Y(N28351) );
  OAI222XL U12612 ( .A0(n7436), .A1(n3010), .B0(n3046), .B1(n8088), .C0(n7533), 
        .C1(n8085), .Y(N28415) );
  OAI222XL U12613 ( .A0(n7436), .A1(n8154), .B0(n2563), .B1(n8153), .C0(n7533), 
        .C1(n8149), .Y(N28735) );
  OAI222XL U12614 ( .A0(n7436), .A1(n8167), .B0(n8166), .B1(n2431), .C0(n8163), 
        .C1(n7533), .Y(N28799) );
  OAI222XL U12615 ( .A0(n7438), .A1(n8014), .B0(n3466), .B1(n8011), .C0(n7532), 
        .C1(n8008), .Y(N28032) );
  OAI222XL U12616 ( .A0(n7438), .A1(n3362), .B0(n3397), .B1(n8024), .C0(n7532), 
        .C1(n6612), .Y(N28096) );
  OAI222XL U12617 ( .A0(n7438), .A1(n8078), .B0(n3116), .B1(n8076), .C0(n7532), 
        .C1(n6614), .Y(N28352) );
  OAI222XL U12618 ( .A0(n7438), .A1(n3010), .B0(n3045), .B1(n8088), .C0(n7532), 
        .C1(n8085), .Y(N28416) );
  AOI221XL U12619 ( .A0(n8609), .A1(n8160), .B0(n8610), .B1(n8146), .C0(n4275), 
        .Y(n4263) );
  OAI222XL U12620 ( .A0(n8082), .A1(n3045), .B0(n8018), .B1(n3397), .C0(n8069), 
        .C1(n3116), .Y(n4275) );
  OAI222XL U12621 ( .A0(n8623), .A1(n7934), .B0(n7931), .B1(n9168), .C0(n8005), 
        .C1(n3469), .Y(n4326) );
  OAI222XL U12622 ( .A0(n8618), .A1(n7934), .B0(n7931), .B1(n9160), .C0(n8006), 
        .C1(n3468), .Y(n4308) );
  OAI222XL U12623 ( .A0(n8613), .A1(n7934), .B0(n7931), .B1(n9152), .C0(n3498), 
        .C1(n3467), .Y(n4290) );
  OAI221XL U12624 ( .A0(n7434), .A1(n7990), .B0(n7534), .B1(n7985), .C0(n3606), 
        .Y(N27902) );
  OAI221XL U12625 ( .A0(n7434), .A1(n8054), .B0(n7534), .B1(n8051), .C0(n3260), 
        .Y(N28222) );
  OAI221XL U12626 ( .A0(n7434), .A1(n8105), .B0(n7534), .B1(n8102), .C0(n2977), 
        .Y(N28478) );
  OAI221XL U12627 ( .A0(n7434), .A1(n8118), .B0(n7534), .B1(n8113), .C0(n2875), 
        .Y(N28542) );
  OAI221XL U12628 ( .A0(n7434), .A1(n8131), .B0(n7534), .B1(n8128), .C0(n2770), 
        .Y(N28606) );
  OAI221XL U12629 ( .A0(n7434), .A1(n7977), .B0(n7534), .B1(n7974), .C0(n4297), 
        .Y(N27838) );
  OAI221XL U12630 ( .A0(n7436), .A1(n7988), .B0(n7533), .B1(n7985), .C0(n3605), 
        .Y(N27903) );
  OAI221XL U12631 ( .A0(n7436), .A1(n8054), .B0(n7533), .B1(n8051), .C0(n3259), 
        .Y(N28223) );
  OAI221XL U12632 ( .A0(n7436), .A1(n8105), .B0(n7533), .B1(n8102), .C0(n2976), 
        .Y(N28479) );
  OAI221XL U12633 ( .A0(n7436), .A1(n8118), .B0(n7533), .B1(n8115), .C0(n2873), 
        .Y(N28543) );
  OAI221XL U12634 ( .A0(n7436), .A1(n8131), .B0(n7533), .B1(n8128), .C0(n2769), 
        .Y(N28607) );
  OAI221XL U12635 ( .A0(n7436), .A1(n7977), .B0(n7533), .B1(n7974), .C0(n4279), 
        .Y(N27839) );
  OAI221XL U12636 ( .A0(n7438), .A1(n7988), .B0(n7532), .B1(n7986), .C0(n3604), 
        .Y(N27904) );
  AOI2BB2X1 U12637 ( .B0(n7984), .B1(n7437), .A0N(n9150), .A1N(n7980), .Y(
        n3604) );
  OAI221XL U12638 ( .A0(n7438), .A1(n8054), .B0(n7532), .B1(n8049), .C0(n3258), 
        .Y(N28224) );
  AOI2BB2X1 U12639 ( .B0(n8048), .B1(n7437), .A0N(n9148), .A1N(n8044), .Y(
        n3258) );
  OAI221XL U12640 ( .A0(n7438), .A1(n8103), .B0(n7532), .B1(n8102), .C0(n2975), 
        .Y(N28480) );
  AOI2BB2X1 U12641 ( .B0(n8096), .B1(n7437), .A0N(n9146), .A1N(n8095), .Y(
        n2975) );
  OAI221XL U12642 ( .A0(n7438), .A1(n8118), .B0(n7532), .B1(n8115), .C0(n2871), 
        .Y(N28544) );
  AOI2BB2X1 U12643 ( .B0(n8110), .B1(n7437), .A0N(n9145), .A1N(n8108), .Y(
        n2871) );
  OAI221XL U12644 ( .A0(n7438), .A1(n8129), .B0(n7532), .B1(n8128), .C0(n2768), 
        .Y(N28608) );
  OAI221XL U12645 ( .A0(n7438), .A1(n7977), .B0(n7532), .B1(n7972), .C0(n4261), 
        .Y(N27840) );
  AOI2BB2X1 U12646 ( .B0(n7970), .B1(n7437), .A0N(n9143), .A1N(n7968), .Y(
        n4261) );
  OAI222XL U12647 ( .A0(n9202), .A1(n7941), .B0(n8643), .B1(n7940), .C0(n7937), 
        .C1(n9201), .Y(n4395) );
  OAI222XL U12648 ( .A0(n7958), .A1(n9199), .B0(n9206), .B1(n7954), .C0(n8643), 
        .C1(n7952), .Y(n4393) );
  OAI222XL U12649 ( .A0(n9194), .A1(n7942), .B0(n8638), .B1(n7940), .C0(n7937), 
        .C1(n9193), .Y(n4377) );
  OAI222XL U12650 ( .A0(n7957), .A1(n9191), .B0(n9198), .B1(n7955), .C0(n8638), 
        .C1(n7952), .Y(n4375) );
  OAI222XL U12651 ( .A0(n9186), .A1(n7941), .B0(n8633), .B1(n6604), .C0(n7937), 
        .C1(n9185), .Y(n4359) );
  OAI222XL U12652 ( .A0(n7957), .A1(n9183), .B0(n9190), .B1(n7954), .C0(n8633), 
        .C1(n7952), .Y(n4357) );
  OAI222XL U12653 ( .A0(n9178), .A1(n7942), .B0(n8628), .B1(n6604), .C0(n7937), 
        .C1(n9177), .Y(n4341) );
  OAI222XL U12654 ( .A0(n7957), .A1(n9175), .B0(n9182), .B1(n7955), .C0(n8628), 
        .C1(n7952), .Y(n4339) );
  OAI222XL U12655 ( .A0(n9170), .A1(n7943), .B0(n8623), .B1(n7940), .C0(n7937), 
        .C1(n9169), .Y(n4323) );
  OAI222XL U12656 ( .A0(n7957), .A1(n9167), .B0(n9174), .B1(n7953), .C0(n8623), 
        .C1(n7951), .Y(n4321) );
  OAI222XL U12657 ( .A0(n7424), .A1(n6585), .B0(n3541), .B1(n8000), .C0(n7539), 
        .C1(n7995), .Y(N27961) );
  OAI222XL U12658 ( .A0(n7424), .A1(n8013), .B0(n3473), .B1(n8012), .C0(n7539), 
        .C1(n8007), .Y(N28025) );
  OAI222XL U12659 ( .A0(n7424), .A1(n8027), .B0(n3404), .B1(n8025), .C0(n7539), 
        .C1(n8021), .Y(N28089) );
  OAI222XL U12660 ( .A0(n7424), .A1(n8040), .B0(n3336), .B1(n8036), .C0(n7539), 
        .C1(n8034), .Y(N28153) );
  OAI222XL U12661 ( .A0(n7424), .A1(n8077), .B0(n3123), .B1(n8074), .C0(n7539), 
        .C1(n8072), .Y(N28345) );
  OAI222XL U12662 ( .A0(n7424), .A1(n8091), .B0(n3052), .B1(n8089), .C0(n7539), 
        .C1(n8084), .Y(N28409) );
  OAI222XL U12663 ( .A0(n7424), .A1(n6586), .B0(n2569), .B1(n8152), .C0(n7539), 
        .C1(n8148), .Y(N28729) );
  OAI222XL U12664 ( .A0(n7424), .A1(n8168), .B0(n6580), .B1(n2449), .C0(n8161), 
        .C1(n7539), .Y(N28793) );
  OAI222XL U12665 ( .A0(n7426), .A1(n6585), .B0(n3540), .B1(n7998), .C0(n7538), 
        .C1(n7995), .Y(N27962) );
  OAI222XL U12666 ( .A0(n7426), .A1(n8013), .B0(n3472), .B1(n8012), .C0(n7538), 
        .C1(n8007), .Y(N28026) );
  OAI222XL U12667 ( .A0(n7426), .A1(n8027), .B0(n3403), .B1(n8025), .C0(n7538), 
        .C1(n8021), .Y(N28090) );
  OAI222XL U12668 ( .A0(n7426), .A1(n8040), .B0(n3335), .B1(n8038), .C0(n7538), 
        .C1(n8034), .Y(N28154) );
  OAI222XL U12669 ( .A0(n7426), .A1(n8077), .B0(n3122), .B1(n8076), .C0(n7538), 
        .C1(n8072), .Y(N28346) );
  OAI222XL U12670 ( .A0(n7426), .A1(n8091), .B0(n3051), .B1(n8089), .C0(n7538), 
        .C1(n8084), .Y(N28410) );
  OAI222XL U12671 ( .A0(n7426), .A1(n6586), .B0(n2568), .B1(n8151), .C0(n7538), 
        .C1(n8148), .Y(N28730) );
  OAI222XL U12672 ( .A0(n7426), .A1(n8169), .B0(n8166), .B1(n2446), .C0(n8161), 
        .C1(n7538), .Y(N28794) );
  OAI222XL U12673 ( .A0(n7428), .A1(n6585), .B0(n3539), .B1(n7999), .C0(n7537), 
        .C1(n7995), .Y(N27963) );
  OAI222XL U12674 ( .A0(n7428), .A1(n8013), .B0(n3471), .B1(n8012), .C0(n7537), 
        .C1(n8007), .Y(N28027) );
  OAI222XL U12675 ( .A0(n7428), .A1(n8027), .B0(n3402), .B1(n8025), .C0(n7537), 
        .C1(n8021), .Y(N28091) );
  OAI222XL U12676 ( .A0(n7428), .A1(n8040), .B0(n3334), .B1(n8037), .C0(n7537), 
        .C1(n8034), .Y(N28155) );
  OAI222XL U12677 ( .A0(n7428), .A1(n8077), .B0(n3121), .B1(n8075), .C0(n7537), 
        .C1(n8072), .Y(N28347) );
  OAI222XL U12678 ( .A0(n7428), .A1(n8091), .B0(n3050), .B1(n8089), .C0(n7537), 
        .C1(n8084), .Y(N28411) );
  OAI222XL U12679 ( .A0(n7428), .A1(n6586), .B0(n2567), .B1(n8153), .C0(n7537), 
        .C1(n8148), .Y(N28731) );
  OAI222XL U12680 ( .A0(n7428), .A1(n8169), .B0(n8166), .B1(n2443), .C0(n8161), 
        .C1(n7537), .Y(N28795) );
  OAI222XL U12681 ( .A0(n7430), .A1(n6585), .B0(n3538), .B1(n8000), .C0(n7536), 
        .C1(n7995), .Y(N27964) );
  OAI222XL U12682 ( .A0(n7430), .A1(n8013), .B0(n3470), .B1(n8012), .C0(n7536), 
        .C1(n8007), .Y(N28028) );
  OAI222XL U12683 ( .A0(n7430), .A1(n8027), .B0(n3401), .B1(n8025), .C0(n7536), 
        .C1(n8021), .Y(N28092) );
  OAI222XL U12684 ( .A0(n7430), .A1(n8040), .B0(n3333), .B1(n8036), .C0(n7536), 
        .C1(n8034), .Y(N28156) );
  OAI222XL U12685 ( .A0(n7430), .A1(n8077), .B0(n3120), .B1(n8074), .C0(n7536), 
        .C1(n8072), .Y(N28348) );
  OAI222XL U12686 ( .A0(n7430), .A1(n8091), .B0(n3049), .B1(n8089), .C0(n7536), 
        .C1(n8084), .Y(N28412) );
  OAI222XL U12687 ( .A0(n7430), .A1(n6586), .B0(n2566), .B1(n8152), .C0(n7536), 
        .C1(n8148), .Y(N28732) );
  OAI222XL U12688 ( .A0(n7430), .A1(n8169), .B0(n8166), .B1(n2440), .C0(n8161), 
        .C1(n7536), .Y(N28796) );
  OAI222XL U12689 ( .A0(n8643), .A1(n7934), .B0(n7930), .B1(n9200), .C0(n8005), 
        .C1(n3473), .Y(n4398) );
  OAI222XL U12690 ( .A0(n8638), .A1(n3675), .B0(n7931), .B1(n9192), .C0(n8005), 
        .C1(n3472), .Y(n4380) );
  OAI222XL U12691 ( .A0(n8633), .A1(n3675), .B0(n7931), .B1(n9184), .C0(n3498), 
        .C1(n3471), .Y(n4362) );
  OAI222XL U12692 ( .A0(n8628), .A1(n3675), .B0(n7931), .B1(n9176), .C0(n3498), 
        .C1(n3470), .Y(n4344) );
  OAI221XL U12693 ( .A0(n7424), .A1(n7988), .B0(n7539), .B1(n7986), .C0(n3611), 
        .Y(N27897) );
  OAI221XL U12694 ( .A0(n7424), .A1(n8052), .B0(n7539), .B1(n8050), .C0(n3265), 
        .Y(N28217) );
  OAI221XL U12695 ( .A0(n7424), .A1(n8103), .B0(n7539), .B1(n8100), .C0(n2982), 
        .Y(N28473) );
  OAI221XL U12696 ( .A0(n7424), .A1(n8116), .B0(n7539), .B1(n8113), .C0(n2885), 
        .Y(N28537) );
  OAI221XL U12697 ( .A0(n7424), .A1(n8130), .B0(n7539), .B1(n8126), .C0(n2775), 
        .Y(N28601) );
  OAI221XL U12698 ( .A0(n7424), .A1(n7976), .B0(n7539), .B1(n7973), .C0(n4387), 
        .Y(N27833) );
  OAI221XL U12699 ( .A0(n7426), .A1(n7988), .B0(n7538), .B1(n7986), .C0(n3610), 
        .Y(N27898) );
  OAI221XL U12700 ( .A0(n7426), .A1(n8052), .B0(n7538), .B1(n8051), .C0(n3264), 
        .Y(N28218) );
  OAI221XL U12701 ( .A0(n7426), .A1(n8103), .B0(n7538), .B1(n8102), .C0(n2981), 
        .Y(N28474) );
  OAI221XL U12702 ( .A0(n7426), .A1(n8116), .B0(n7538), .B1(n8115), .C0(n2883), 
        .Y(N28538) );
  OAI221XL U12703 ( .A0(n7426), .A1(n8130), .B0(n7538), .B1(n6600), .C0(n2774), 
        .Y(N28602) );
  OAI221XL U12704 ( .A0(n7426), .A1(n7976), .B0(n7538), .B1(n7972), .C0(n4369), 
        .Y(N27834) );
  OAI221XL U12705 ( .A0(n7428), .A1(n7988), .B0(n7537), .B1(n7987), .C0(n3609), 
        .Y(N27899) );
  OAI221XL U12706 ( .A0(n7428), .A1(n8054), .B0(n7537), .B1(n8051), .C0(n3263), 
        .Y(N28219) );
  OAI221XL U12707 ( .A0(n7428), .A1(n8103), .B0(n7537), .B1(n8102), .C0(n2980), 
        .Y(N28475) );
  OAI221XL U12708 ( .A0(n7428), .A1(n8118), .B0(n7537), .B1(n8115), .C0(n2881), 
        .Y(N28539) );
  OAI221XL U12709 ( .A0(n7428), .A1(n6609), .B0(n7537), .B1(n6600), .C0(n2773), 
        .Y(N28603) );
  OAI221XL U12710 ( .A0(n7428), .A1(n7977), .B0(n7537), .B1(n7972), .C0(n4351), 
        .Y(N27835) );
  OAI221XL U12711 ( .A0(n7430), .A1(n7990), .B0(n7536), .B1(n7985), .C0(n3608), 
        .Y(N27900) );
  OAI221XL U12712 ( .A0(n7430), .A1(n8054), .B0(n7536), .B1(n8049), .C0(n3262), 
        .Y(N28220) );
  OAI221XL U12713 ( .A0(n7430), .A1(n8103), .B0(n7536), .B1(n8102), .C0(n2979), 
        .Y(N28476) );
  OAI221XL U12714 ( .A0(n7430), .A1(n8118), .B0(n7536), .B1(n8115), .C0(n2879), 
        .Y(N28540) );
  OAI221XL U12715 ( .A0(n7430), .A1(n8129), .B0(n7536), .B1(n8128), .C0(n2772), 
        .Y(N28604) );
  OAI221XL U12716 ( .A0(n7430), .A1(n7977), .B0(n7536), .B1(n7972), .C0(n4333), 
        .Y(N27836) );
  OAI221XL U12717 ( .A0(n7432), .A1(n7990), .B0(n7535), .B1(n7985), .C0(n3607), 
        .Y(N27901) );
  OAI221XL U12718 ( .A0(n7432), .A1(n8054), .B0(n7535), .B1(n8051), .C0(n3261), 
        .Y(N28221) );
  OAI221XL U12719 ( .A0(n7432), .A1(n8103), .B0(n7535), .B1(n8102), .C0(n2978), 
        .Y(N28477) );
  OAI221XL U12720 ( .A0(n7432), .A1(n8118), .B0(n7535), .B1(n8115), .C0(n2877), 
        .Y(N28541) );
  OAI221XL U12721 ( .A0(n7432), .A1(n6609), .B0(n7535), .B1(n8126), .C0(n2771), 
        .Y(N28605) );
  OAI221XL U12722 ( .A0(n7432), .A1(n7977), .B0(n7535), .B1(n7972), .C0(n4315), 
        .Y(N27837) );
  OAI222XL U12723 ( .A0(n8658), .A1(n7933), .B0(n7929), .B1(n9224), .C0(n8005), 
        .C1(n3476), .Y(n4452) );
  OAI222XL U12724 ( .A0(n7958), .A1(n9223), .B0(n9230), .B1(n7955), .C0(n8658), 
        .C1(n7952), .Y(n4447) );
  OAI222XL U12725 ( .A0(n8653), .A1(n7933), .B0(n7930), .B1(n9216), .C0(n8005), 
        .C1(n3475), .Y(n4434) );
  OAI222XL U12726 ( .A0(n7958), .A1(n9215), .B0(n9222), .B1(n7955), .C0(n8653), 
        .C1(n7952), .Y(n4429) );
  OAI222XL U12727 ( .A0(n9210), .A1(n7941), .B0(n8648), .B1(n7940), .C0(n7937), 
        .C1(n9209), .Y(n4413) );
  OAI222XL U12728 ( .A0(n7958), .A1(n9207), .B0(n9214), .B1(n7955), .C0(n8648), 
        .C1(n7952), .Y(n4411) );
  OAI222XL U12729 ( .A0(n7418), .A1(n8003), .B0(n3544), .B1(n6581), .C0(n7542), 
        .C1(n7995), .Y(N27958) );
  OAI222XL U12730 ( .A0(n7418), .A1(n8013), .B0(n3476), .B1(n8012), .C0(n7542), 
        .C1(n8007), .Y(N28022) );
  OAI222XL U12731 ( .A0(n7418), .A1(n8027), .B0(n3407), .B1(n8025), .C0(n7542), 
        .C1(n8021), .Y(N28086) );
  OAI222XL U12732 ( .A0(n7418), .A1(n8040), .B0(n3339), .B1(n8038), .C0(n7542), 
        .C1(n8034), .Y(N28150) );
  OAI222XL U12733 ( .A0(n7418), .A1(n8077), .B0(n3126), .B1(n8076), .C0(n7542), 
        .C1(n8072), .Y(N28342) );
  OAI222XL U12734 ( .A0(n7418), .A1(n8091), .B0(n3055), .B1(n8089), .C0(n7542), 
        .C1(n8084), .Y(N28406) );
  OAI222XL U12735 ( .A0(n7418), .A1(n8156), .B0(n2572), .B1(n6587), .C0(n7542), 
        .C1(n8148), .Y(N28726) );
  OAI222XL U12736 ( .A0(n7418), .A1(n8167), .B0(n8166), .B1(n2458), .C0(n8161), 
        .C1(n7542), .Y(N28790) );
  OAI222XL U12737 ( .A0(n7420), .A1(n6585), .B0(n3543), .B1(n7998), .C0(n7541), 
        .C1(n7995), .Y(N27959) );
  OAI222XL U12738 ( .A0(n7420), .A1(n8013), .B0(n3475), .B1(n8012), .C0(n7541), 
        .C1(n8007), .Y(N28023) );
  OAI222XL U12739 ( .A0(n7420), .A1(n8027), .B0(n3406), .B1(n8025), .C0(n7541), 
        .C1(n8021), .Y(N28087) );
  OAI222XL U12740 ( .A0(n7420), .A1(n8040), .B0(n3338), .B1(n8037), .C0(n7541), 
        .C1(n8034), .Y(N28151) );
  OAI222XL U12741 ( .A0(n7420), .A1(n8077), .B0(n3125), .B1(n8075), .C0(n7541), 
        .C1(n8072), .Y(N28343) );
  OAI222XL U12742 ( .A0(n7420), .A1(n8091), .B0(n3054), .B1(n8089), .C0(n7541), 
        .C1(n8084), .Y(N28407) );
  OAI222XL U12743 ( .A0(n7420), .A1(n6586), .B0(n2571), .B1(n8151), .C0(n7541), 
        .C1(n8148), .Y(N28727) );
  OAI222XL U12744 ( .A0(n7420), .A1(n6588), .B0(n6580), .B1(n2455), .C0(n8161), 
        .C1(n7541), .Y(N28791) );
  OAI222XL U12745 ( .A0(n7422), .A1(n6585), .B0(n3542), .B1(n7999), .C0(n7540), 
        .C1(n7995), .Y(N27960) );
  OAI222XL U12746 ( .A0(n7422), .A1(n8013), .B0(n3474), .B1(n8012), .C0(n7540), 
        .C1(n8007), .Y(N28024) );
  OAI222XL U12747 ( .A0(n7422), .A1(n8027), .B0(n3405), .B1(n8025), .C0(n7540), 
        .C1(n8021), .Y(N28088) );
  OAI222XL U12748 ( .A0(n7422), .A1(n8040), .B0(n3337), .B1(n8036), .C0(n7540), 
        .C1(n8034), .Y(N28152) );
  OAI222XL U12749 ( .A0(n7422), .A1(n8077), .B0(n3124), .B1(n8074), .C0(n7540), 
        .C1(n8072), .Y(N28344) );
  OAI222XL U12750 ( .A0(n7422), .A1(n8091), .B0(n3053), .B1(n8089), .C0(n7540), 
        .C1(n8084), .Y(N28408) );
  OAI222XL U12751 ( .A0(n7422), .A1(n6586), .B0(n2570), .B1(n8153), .C0(n7540), 
        .C1(n8148), .Y(N28728) );
  OAI222XL U12752 ( .A0(n7422), .A1(n6588), .B0(n6580), .B1(n2452), .C0(n8161), 
        .C1(n7540), .Y(N28792) );
  AOI221XL U12753 ( .A0(n8659), .A1(n8157), .B0(n8660), .B1(n8145), .C0(n4455), 
        .Y(n4443) );
  CLKINVX1 U12754 ( .A(n2458), .Y(n8659) );
  CLKINVX1 U12755 ( .A(n2572), .Y(n8660) );
  OAI222XL U12756 ( .A0(n8081), .A1(n3055), .B0(n8017), .B1(n3407), .C0(n8069), 
        .C1(n3126), .Y(n4455) );
  AOI221XL U12757 ( .A0(n8654), .A1(n6610), .B0(n8655), .B1(n8145), .C0(n4437), 
        .Y(n4425) );
  CLKINVX1 U12758 ( .A(n2455), .Y(n8654) );
  CLKINVX1 U12759 ( .A(n2571), .Y(n8655) );
  OAI222XL U12760 ( .A0(n8081), .A1(n3054), .B0(n8017), .B1(n3406), .C0(n8069), 
        .C1(n3125), .Y(n4437) );
  CLKINVX1 U12761 ( .A(n2452), .Y(n8649) );
  CLKINVX1 U12762 ( .A(n2570), .Y(n8650) );
  CLKINVX1 U12763 ( .A(n3542), .Y(n8651) );
  CLKINVX1 U12764 ( .A(n3337), .Y(n8652) );
  OAI222XL U12765 ( .A0(n8648), .A1(n7932), .B0(n7930), .B1(n9208), .C0(n8005), 
        .C1(n3474), .Y(n4416) );
  OAI221XL U12766 ( .A0(n7418), .A1(n7988), .B0(n7542), .B1(n7985), .C0(n3614), 
        .Y(N27894) );
  OAI221XL U12767 ( .A0(n7418), .A1(n8052), .B0(n7542), .B1(n8050), .C0(n3268), 
        .Y(N28214) );
  OAI221XL U12768 ( .A0(n7418), .A1(n8103), .B0(n7542), .B1(n8100), .C0(n2985), 
        .Y(N28470) );
  OAI221XL U12769 ( .A0(n7418), .A1(n8116), .B0(n7542), .B1(n8113), .C0(n2891), 
        .Y(N28534) );
  OAI221XL U12770 ( .A0(n7418), .A1(n8130), .B0(n7542), .B1(n8126), .C0(n2778), 
        .Y(N28598) );
  OAI221XL U12771 ( .A0(n7418), .A1(n7976), .B0(n7542), .B1(n7972), .C0(n4441), 
        .Y(N27830) );
  OAI221XL U12772 ( .A0(n7420), .A1(n7988), .B0(n7541), .B1(n7986), .C0(n3613), 
        .Y(N27895) );
  OAI221XL U12773 ( .A0(n7420), .A1(n8052), .B0(n7541), .B1(n8050), .C0(n3267), 
        .Y(N28215) );
  OAI221XL U12774 ( .A0(n7420), .A1(n8103), .B0(n7541), .B1(n8100), .C0(n2984), 
        .Y(N28471) );
  OAI221XL U12775 ( .A0(n7420), .A1(n8116), .B0(n7541), .B1(n8113), .C0(n2889), 
        .Y(N28535) );
  OAI221XL U12776 ( .A0(n7420), .A1(n8130), .B0(n7541), .B1(n8126), .C0(n2777), 
        .Y(N28599) );
  OAI221XL U12777 ( .A0(n7420), .A1(n7976), .B0(n7541), .B1(n7973), .C0(n4423), 
        .Y(N27831) );
  OAI221XL U12778 ( .A0(n7422), .A1(n7988), .B0(n7540), .B1(n7986), .C0(n3612), 
        .Y(N27896) );
  OAI221XL U12779 ( .A0(n7422), .A1(n8052), .B0(n7540), .B1(n8050), .C0(n3266), 
        .Y(N28216) );
  OAI221XL U12780 ( .A0(n7422), .A1(n8103), .B0(n7540), .B1(n8100), .C0(n2983), 
        .Y(N28472) );
  OAI221XL U12781 ( .A0(n7422), .A1(n8116), .B0(n7540), .B1(n8113), .C0(n2887), 
        .Y(N28536) );
  OAI221XL U12782 ( .A0(n7422), .A1(n8130), .B0(n7540), .B1(n8126), .C0(n2776), 
        .Y(N28600) );
  OAI221XL U12783 ( .A0(n7422), .A1(n7976), .B0(n7540), .B1(n7973), .C0(n4405), 
        .Y(N27832) );
  CLKINVX1 U12784 ( .A(n3339), .Y(n8662) );
  CLKINVX1 U12785 ( .A(n3338), .Y(n8657) );
  CLKINVX1 U12786 ( .A(n3544), .Y(n8661) );
  CLKINVX1 U12787 ( .A(n3543), .Y(n8656) );
  OAI222XL U12788 ( .A0(n9266), .A1(n7941), .B0(n8683), .B1(n7938), .C0(n7937), 
        .C1(n9265), .Y(n4539) );
  OAI222XL U12789 ( .A0(n7958), .A1(n9263), .B0(n9270), .B1(n7955), .C0(n8683), 
        .C1(n7952), .Y(n4537) );
  OAI222XL U12790 ( .A0(n9258), .A1(n7942), .B0(n8678), .B1(n7940), .C0(n3671), 
        .C1(n9257), .Y(n4521) );
  OAI222XL U12791 ( .A0(n7958), .A1(n9255), .B0(n9262), .B1(n7953), .C0(n8678), 
        .C1(n7952), .Y(n4519) );
  OAI222XL U12792 ( .A0(n9250), .A1(n7941), .B0(n8673), .B1(n7938), .C0(n3671), 
        .C1(n9249), .Y(n4503) );
  OAI222XL U12793 ( .A0(n7958), .A1(n9247), .B0(n9254), .B1(n7954), .C0(n8673), 
        .C1(n7952), .Y(n4501) );
  OAI222XL U12794 ( .A0(n9242), .A1(n7942), .B0(n8668), .B1(n7939), .C0(n3671), 
        .C1(n9241), .Y(n4485) );
  OAI222XL U12795 ( .A0(n7958), .A1(n9239), .B0(n9246), .B1(n7955), .C0(n8668), 
        .C1(n7952), .Y(n4483) );
  OAI222XL U12796 ( .A0(n9234), .A1(n7941), .B0(n8663), .B1(n7939), .C0(n7937), 
        .C1(n9233), .Y(n4467) );
  OAI222XL U12797 ( .A0(n7958), .A1(n9231), .B0(n9238), .B1(n7954), .C0(n8663), 
        .C1(n7952), .Y(n4465) );
  OAI222XL U12798 ( .A0(n7406), .A1(n8003), .B0(n3550), .B1(n7999), .C0(n7548), 
        .C1(n7995), .Y(N27952) );
  OAI222XL U12799 ( .A0(n7406), .A1(n8013), .B0(n3482), .B1(n8012), .C0(n7548), 
        .C1(n8007), .Y(N28016) );
  OAI222XL U12800 ( .A0(n7406), .A1(n8027), .B0(n3413), .B1(n8025), .C0(n7548), 
        .C1(n8021), .Y(N28080) );
  OAI222XL U12801 ( .A0(n7406), .A1(n8040), .B0(n3345), .B1(n8037), .C0(n7548), 
        .C1(n8034), .Y(N28144) );
  OAI222XL U12802 ( .A0(n7406), .A1(n8077), .B0(n3132), .B1(n8075), .C0(n7548), 
        .C1(n8072), .Y(N28336) );
  OAI222XL U12803 ( .A0(n7406), .A1(n8091), .B0(n3061), .B1(n8087), .C0(n7548), 
        .C1(n8084), .Y(N28400) );
  OAI222XL U12804 ( .A0(n7406), .A1(n8156), .B0(n2578), .B1(n8152), .C0(n7548), 
        .C1(n8148), .Y(N28720) );
  OAI222XL U12805 ( .A0(n7406), .A1(n6588), .B0(n6580), .B1(n2476), .C0(n8161), 
        .C1(n7548), .Y(N28784) );
  OAI222XL U12806 ( .A0(n7408), .A1(n8002), .B0(n3549), .B1(n7998), .C0(n7547), 
        .C1(n7995), .Y(N27953) );
  OAI222XL U12807 ( .A0(n7408), .A1(n8013), .B0(n3481), .B1(n8012), .C0(n7547), 
        .C1(n8007), .Y(N28017) );
  OAI222XL U12808 ( .A0(n7408), .A1(n8027), .B0(n3412), .B1(n8025), .C0(n7547), 
        .C1(n8021), .Y(N28081) );
  OAI222XL U12809 ( .A0(n7408), .A1(n8040), .B0(n3344), .B1(n8037), .C0(n7547), 
        .C1(n8034), .Y(N28145) );
  OAI222XL U12810 ( .A0(n7408), .A1(n8077), .B0(n3131), .B1(n8075), .C0(n7547), 
        .C1(n8072), .Y(N28337) );
  OAI222XL U12811 ( .A0(n7408), .A1(n8091), .B0(n3060), .B1(n8089), .C0(n7547), 
        .C1(n8084), .Y(N28401) );
  OAI222XL U12812 ( .A0(n7408), .A1(n8155), .B0(n2577), .B1(n8152), .C0(n7547), 
        .C1(n8148), .Y(N28721) );
  OAI222XL U12813 ( .A0(n7408), .A1(n6588), .B0(n6580), .B1(n2473), .C0(n8161), 
        .C1(n7547), .Y(N28785) );
  OAI222XL U12814 ( .A0(n7410), .A1(n8003), .B0(n3548), .B1(n7999), .C0(n7546), 
        .C1(n7995), .Y(N27954) );
  OAI222XL U12815 ( .A0(n7410), .A1(n8013), .B0(n3480), .B1(n8012), .C0(n7546), 
        .C1(n8007), .Y(N28018) );
  OAI222XL U12816 ( .A0(n7410), .A1(n8027), .B0(n3411), .B1(n8025), .C0(n7546), 
        .C1(n8021), .Y(N28082) );
  OAI222XL U12817 ( .A0(n7410), .A1(n8040), .B0(n3343), .B1(n8036), .C0(n7546), 
        .C1(n8034), .Y(N28146) );
  OAI222XL U12818 ( .A0(n7410), .A1(n8077), .B0(n3130), .B1(n8074), .C0(n7546), 
        .C1(n8072), .Y(N28338) );
  OAI222XL U12819 ( .A0(n7410), .A1(n8091), .B0(n3059), .B1(n8089), .C0(n7546), 
        .C1(n8084), .Y(N28402) );
  OAI222XL U12820 ( .A0(n7410), .A1(n8156), .B0(n2576), .B1(n8151), .C0(n7546), 
        .C1(n8148), .Y(N28722) );
  OAI222XL U12821 ( .A0(n7410), .A1(n8168), .B0(n8164), .B1(n2470), .C0(n8161), 
        .C1(n7546), .Y(N28786) );
  OAI222XL U12822 ( .A0(n7412), .A1(n8002), .B0(n3547), .B1(n8000), .C0(n7545), 
        .C1(n7995), .Y(N27955) );
  OAI222XL U12823 ( .A0(n7412), .A1(n8013), .B0(n3479), .B1(n8012), .C0(n7545), 
        .C1(n8007), .Y(N28019) );
  OAI222XL U12824 ( .A0(n7412), .A1(n8027), .B0(n3410), .B1(n8025), .C0(n7545), 
        .C1(n8021), .Y(N28083) );
  OAI222XL U12825 ( .A0(n7412), .A1(n8040), .B0(n3342), .B1(n6575), .C0(n7545), 
        .C1(n8034), .Y(N28147) );
  OAI222XL U12826 ( .A0(n7412), .A1(n8077), .B0(n3129), .B1(n6590), .C0(n7545), 
        .C1(n8072), .Y(N28339) );
  OAI222XL U12827 ( .A0(n7412), .A1(n8091), .B0(n3058), .B1(n8089), .C0(n7545), 
        .C1(n8084), .Y(N28403) );
  OAI222XL U12828 ( .A0(n7412), .A1(n8155), .B0(n2575), .B1(n8153), .C0(n7545), 
        .C1(n8148), .Y(N28723) );
  OAI222XL U12829 ( .A0(n7412), .A1(n8167), .B0(n8164), .B1(n2467), .C0(n8161), 
        .C1(n7545), .Y(N28787) );
  OAI222XL U12830 ( .A0(n7414), .A1(n8003), .B0(n3546), .B1(n7998), .C0(n7544), 
        .C1(n7995), .Y(N27956) );
  OAI222XL U12831 ( .A0(n7414), .A1(n8013), .B0(n3478), .B1(n8012), .C0(n7544), 
        .C1(n8007), .Y(N28020) );
  OAI222XL U12832 ( .A0(n7414), .A1(n8027), .B0(n3409), .B1(n8025), .C0(n7544), 
        .C1(n8021), .Y(N28084) );
  OAI222XL U12833 ( .A0(n7414), .A1(n8040), .B0(n3341), .B1(n8038), .C0(n7544), 
        .C1(n8034), .Y(N28148) );
  OAI222XL U12834 ( .A0(n7414), .A1(n8077), .B0(n3128), .B1(n8076), .C0(n7544), 
        .C1(n8072), .Y(N28340) );
  OAI222XL U12835 ( .A0(n7414), .A1(n8091), .B0(n3057), .B1(n8089), .C0(n7544), 
        .C1(n8084), .Y(N28404) );
  OAI222XL U12836 ( .A0(n7414), .A1(n8156), .B0(n2574), .B1(n6587), .C0(n7544), 
        .C1(n8148), .Y(N28724) );
  OAI222XL U12837 ( .A0(n7414), .A1(n8167), .B0(n8165), .B1(n2464), .C0(n8161), 
        .C1(n7544), .Y(N28788) );
  OAI222XL U12838 ( .A0(n7416), .A1(n8002), .B0(n3545), .B1(n7999), .C0(n7543), 
        .C1(n7995), .Y(N27957) );
  OAI222XL U12839 ( .A0(n7416), .A1(n8013), .B0(n3477), .B1(n8012), .C0(n7543), 
        .C1(n8007), .Y(N28021) );
  OAI222XL U12840 ( .A0(n7416), .A1(n8027), .B0(n3408), .B1(n8025), .C0(n7543), 
        .C1(n8021), .Y(N28085) );
  OAI222XL U12841 ( .A0(n7416), .A1(n8040), .B0(n3340), .B1(n8037), .C0(n7543), 
        .C1(n8034), .Y(N28149) );
  OAI222XL U12842 ( .A0(n7416), .A1(n8077), .B0(n3127), .B1(n8075), .C0(n7543), 
        .C1(n8072), .Y(N28341) );
  OAI222XL U12843 ( .A0(n7416), .A1(n8091), .B0(n3056), .B1(n8089), .C0(n7543), 
        .C1(n8084), .Y(N28405) );
  OAI222XL U12844 ( .A0(n7416), .A1(n8155), .B0(n2573), .B1(n6587), .C0(n7543), 
        .C1(n8148), .Y(N28725) );
  OAI222XL U12845 ( .A0(n7416), .A1(n8168), .B0(n8164), .B1(n2461), .C0(n8161), 
        .C1(n7543), .Y(N28789) );
  AOI221XL U12846 ( .A0(n8689), .A1(n8158), .B0(n8690), .B1(n8145), .C0(n4563), 
        .Y(n4551) );
  CLKINVX1 U12847 ( .A(n2476), .Y(n8689) );
  CLKINVX1 U12848 ( .A(n2578), .Y(n8690) );
  OAI222XL U12849 ( .A0(n8081), .A1(n3061), .B0(n8017), .B1(n3413), .C0(n8069), 
        .C1(n3132), .Y(n4563) );
  AOI221XL U12850 ( .A0(n8684), .A1(n6610), .B0(n8685), .B1(n8145), .C0(n4545), 
        .Y(n4533) );
  CLKINVX1 U12851 ( .A(n2473), .Y(n8684) );
  CLKINVX1 U12852 ( .A(n2577), .Y(n8685) );
  OAI222XL U12853 ( .A0(n8081), .A1(n3060), .B0(n8017), .B1(n3412), .C0(n8067), 
        .C1(n3131), .Y(n4545) );
  AOI221XL U12854 ( .A0(n8679), .A1(n8157), .B0(n8680), .B1(n8145), .C0(n4527), 
        .Y(n4515) );
  CLKINVX1 U12855 ( .A(n2470), .Y(n8679) );
  CLKINVX1 U12856 ( .A(n2576), .Y(n8680) );
  OAI222XL U12857 ( .A0(n8081), .A1(n3059), .B0(n8017), .B1(n3411), .C0(n8067), 
        .C1(n3130), .Y(n4527) );
  AOI221XL U12858 ( .A0(n8674), .A1(n8157), .B0(n8675), .B1(n8145), .C0(n4509), 
        .Y(n4497) );
  CLKINVX1 U12859 ( .A(n2467), .Y(n8674) );
  CLKINVX1 U12860 ( .A(n2575), .Y(n8675) );
  OAI222XL U12861 ( .A0(n8081), .A1(n3058), .B0(n8017), .B1(n3410), .C0(n8067), 
        .C1(n3129), .Y(n4509) );
  AOI221XL U12862 ( .A0(n8669), .A1(n8157), .B0(n8670), .B1(n8145), .C0(n4491), 
        .Y(n4479) );
  CLKINVX1 U12863 ( .A(n2464), .Y(n8669) );
  CLKINVX1 U12864 ( .A(n2574), .Y(n8670) );
  OAI222XL U12865 ( .A0(n8081), .A1(n3057), .B0(n8017), .B1(n3409), .C0(n3149), 
        .C1(n3128), .Y(n4491) );
  AOI221XL U12866 ( .A0(n8664), .A1(n8157), .B0(n8665), .B1(n8145), .C0(n4473), 
        .Y(n4461) );
  CLKINVX1 U12867 ( .A(n2461), .Y(n8664) );
  CLKINVX1 U12868 ( .A(n2573), .Y(n8665) );
  OAI222XL U12869 ( .A0(n8081), .A1(n3056), .B0(n8017), .B1(n3408), .C0(n8069), 
        .C1(n3127), .Y(n4473) );
  CLKINVX1 U12870 ( .A(n3549), .Y(n8686) );
  CLKINVX1 U12871 ( .A(n3344), .Y(n8687) );
  OAI222XL U12872 ( .A0(n8683), .A1(n7932), .B0(n3676), .B1(n9264), .C0(n8005), 
        .C1(n3481), .Y(n4542) );
  CLKINVX1 U12873 ( .A(n3548), .Y(n8681) );
  CLKINVX1 U12874 ( .A(n3343), .Y(n8682) );
  OAI222XL U12875 ( .A0(n8678), .A1(n7933), .B0(n7931), .B1(n9256), .C0(n8005), 
        .C1(n3480), .Y(n4524) );
  AOI221XL U12876 ( .A0(n8676), .A1(n7993), .B0(n8677), .B1(n8030), .C0(n4506), 
        .Y(n4498) );
  CLKINVX1 U12877 ( .A(n3547), .Y(n8676) );
  CLKINVX1 U12878 ( .A(n3342), .Y(n8677) );
  OAI222XL U12879 ( .A0(n8673), .A1(n7932), .B0(n7929), .B1(n9248), .C0(n8005), 
        .C1(n3479), .Y(n4506) );
  AOI221XL U12880 ( .A0(n8671), .A1(n7993), .B0(n8672), .B1(n8030), .C0(n4488), 
        .Y(n4480) );
  CLKINVX1 U12881 ( .A(n3546), .Y(n8671) );
  CLKINVX1 U12882 ( .A(n3341), .Y(n8672) );
  OAI222XL U12883 ( .A0(n8668), .A1(n7934), .B0(n7929), .B1(n9240), .C0(n8005), 
        .C1(n3478), .Y(n4488) );
  AOI221XL U12884 ( .A0(n8666), .A1(n7993), .B0(n8667), .B1(n8030), .C0(n4470), 
        .Y(n4462) );
  CLKINVX1 U12885 ( .A(n3545), .Y(n8666) );
  CLKINVX1 U12886 ( .A(n3340), .Y(n8667) );
  OAI222XL U12887 ( .A0(n8663), .A1(n7933), .B0(n7929), .B1(n9232), .C0(n8005), 
        .C1(n3477), .Y(n4470) );
  OAI221XL U12888 ( .A0(n7408), .A1(n6584), .B0(n7547), .B1(n7985), .C0(n3619), 
        .Y(N27889) );
  OAI221XL U12889 ( .A0(n7408), .A1(n6583), .B0(n7547), .B1(n8049), .C0(n3273), 
        .Y(N28209) );
  OAI221XL U12890 ( .A0(n7408), .A1(n8103), .B0(n7547), .B1(n8100), .C0(n2990), 
        .Y(N28465) );
  OAI221XL U12891 ( .A0(n7408), .A1(n8116), .B0(n7547), .B1(n8113), .C0(n2901), 
        .Y(N28529) );
  OAI221XL U12892 ( .A0(n7408), .A1(n8130), .B0(n7547), .B1(n8126), .C0(n2783), 
        .Y(N28593) );
  OAI221XL U12893 ( .A0(n7408), .A1(n7976), .B0(n7547), .B1(n7972), .C0(n4531), 
        .Y(N27825) );
  OAI221XL U12894 ( .A0(n7410), .A1(n6584), .B0(n7546), .B1(n7985), .C0(n3618), 
        .Y(N27890) );
  OAI221XL U12895 ( .A0(n7410), .A1(n6583), .B0(n7546), .B1(n8049), .C0(n3272), 
        .Y(N28210) );
  OAI221XL U12896 ( .A0(n7410), .A1(n6605), .B0(n7546), .B1(n8100), .C0(n2989), 
        .Y(N28466) );
  OAI221XL U12897 ( .A0(n7410), .A1(n6606), .B0(n7546), .B1(n8113), .C0(n2899), 
        .Y(N28530) );
  OAI221XL U12898 ( .A0(n7410), .A1(n8130), .B0(n7546), .B1(n8126), .C0(n2782), 
        .Y(N28594) );
  OAI221XL U12899 ( .A0(n7410), .A1(n7976), .B0(n7546), .B1(n7972), .C0(n4513), 
        .Y(N27826) );
  OAI221XL U12900 ( .A0(n7412), .A1(n6584), .B0(n7545), .B1(n7985), .C0(n3617), 
        .Y(N27891) );
  OAI221XL U12901 ( .A0(n7412), .A1(n6583), .B0(n7545), .B1(n8049), .C0(n3271), 
        .Y(N28211) );
  OAI221XL U12902 ( .A0(n7412), .A1(n6605), .B0(n7545), .B1(n8100), .C0(n2988), 
        .Y(N28467) );
  OAI221XL U12903 ( .A0(n7412), .A1(n6606), .B0(n7545), .B1(n8113), .C0(n2897), 
        .Y(N28531) );
  OAI221XL U12904 ( .A0(n7412), .A1(n8130), .B0(n7545), .B1(n8126), .C0(n2781), 
        .Y(N28595) );
  OAI221XL U12905 ( .A0(n7412), .A1(n7976), .B0(n7545), .B1(n7972), .C0(n4495), 
        .Y(N27827) );
  OAI221XL U12906 ( .A0(n7414), .A1(n6584), .B0(n7544), .B1(n7985), .C0(n3616), 
        .Y(N27892) );
  OAI221XL U12907 ( .A0(n7414), .A1(n6583), .B0(n7544), .B1(n8049), .C0(n3270), 
        .Y(N28212) );
  OAI221XL U12908 ( .A0(n7414), .A1(n6605), .B0(n7544), .B1(n8100), .C0(n2987), 
        .Y(N28468) );
  OAI221XL U12909 ( .A0(n7414), .A1(n6606), .B0(n7544), .B1(n8113), .C0(n2895), 
        .Y(N28532) );
  OAI221XL U12910 ( .A0(n7414), .A1(n8130), .B0(n7544), .B1(n8126), .C0(n2780), 
        .Y(N28596) );
  OAI221XL U12911 ( .A0(n7414), .A1(n7976), .B0(n7544), .B1(n7972), .C0(n4477), 
        .Y(N27828) );
  OAI221XL U12912 ( .A0(n7416), .A1(n6584), .B0(n7543), .B1(n7985), .C0(n3615), 
        .Y(N27893) );
  OAI221XL U12913 ( .A0(n7416), .A1(n8052), .B0(n7543), .B1(n8049), .C0(n3269), 
        .Y(N28213) );
  OAI221XL U12914 ( .A0(n7416), .A1(n8103), .B0(n7543), .B1(n8100), .C0(n2986), 
        .Y(N28469) );
  OAI221XL U12915 ( .A0(n7416), .A1(n6606), .B0(n7543), .B1(n8113), .C0(n2893), 
        .Y(N28533) );
  OAI221XL U12916 ( .A0(n7416), .A1(n8130), .B0(n7543), .B1(n8126), .C0(n2779), 
        .Y(N28597) );
  OAI221XL U12917 ( .A0(n7416), .A1(n7976), .B0(n7543), .B1(n7972), .C0(n4459), 
        .Y(N27829) );
  CLKBUFX3 U12918 ( .A(n6989), .Y(n6977) );
  CLKBUFX3 U12919 ( .A(n8414), .Y(n6989) );
  OAI222XL U12920 ( .A0(n8703), .A1(n7933), .B0(n3676), .B1(n9296), .C0(n8004), 
        .C1(n3485), .Y(n4614) );
  OAI222XL U12921 ( .A0(n7958), .A1(n9295), .B0(n9302), .B1(n7954), .C0(n8703), 
        .C1(n3665), .Y(n4609) );
  OAI222XL U12922 ( .A0(n9290), .A1(n7943), .B0(n8698), .B1(n7939), .C0(n7935), 
        .C1(n9289), .Y(n4593) );
  OAI222XL U12923 ( .A0(n7958), .A1(n9287), .B0(n9294), .B1(n7954), .C0(n8698), 
        .C1(n3665), .Y(n4591) );
  OAI222XL U12924 ( .A0(n9282), .A1(n7943), .B0(n8693), .B1(n7938), .C0(n7937), 
        .C1(n9281), .Y(n4575) );
  OAI222XL U12925 ( .A0(n7958), .A1(n9279), .B0(n9286), .B1(n7954), .C0(n8693), 
        .C1(n7951), .Y(n4573) );
  OAI222XL U12926 ( .A0(n9274), .A1(n7943), .B0(n8688), .B1(n7940), .C0(n7937), 
        .C1(n9273), .Y(n4557) );
  OAI222XL U12927 ( .A0(n7958), .A1(n9271), .B0(n9278), .B1(n7954), .C0(n8688), 
        .C1(n3665), .Y(n4555) );
  OAI222XL U12928 ( .A0(n7400), .A1(n8001), .B0(n3553), .B1(n7998), .C0(n7551), 
        .C1(n6617), .Y(N27949) );
  OAI222XL U12929 ( .A0(n7400), .A1(n3431), .B0(n3485), .B1(n8012), .C0(n7551), 
        .C1(n6618), .Y(N28013) );
  OAI222XL U12930 ( .A0(n7400), .A1(n8026), .B0(n3416), .B1(n8025), .C0(n7551), 
        .C1(n8020), .Y(N28077) );
  OAI222XL U12931 ( .A0(n7400), .A1(n8039), .B0(n3348), .B1(n8036), .C0(n7551), 
        .C1(n8033), .Y(N28141) );
  OAI222XL U12932 ( .A0(n7400), .A1(n3081), .B0(n3135), .B1(n8075), .C0(n7551), 
        .C1(n8071), .Y(N28333) );
  OAI222XL U12933 ( .A0(n7400), .A1(n8090), .B0(n3064), .B1(n8089), .C0(n7551), 
        .C1(n6619), .Y(N28397) );
  OAI222XL U12934 ( .A0(n7400), .A1(n8154), .B0(n2581), .B1(n8151), .C0(n7551), 
        .C1(n6615), .Y(N28717) );
  OAI222XL U12935 ( .A0(n7400), .A1(n8169), .B0(n8164), .B1(n2485), .C0(n8162), 
        .C1(n7551), .Y(N28781) );
  OAI222XL U12936 ( .A0(n7402), .A1(n8003), .B0(n3552), .B1(n8000), .C0(n7550), 
        .C1(n7995), .Y(N27950) );
  OAI222XL U12937 ( .A0(n7402), .A1(n8013), .B0(n3484), .B1(n8010), .C0(n7550), 
        .C1(n8007), .Y(N28014) );
  OAI222XL U12938 ( .A0(n7402), .A1(n8027), .B0(n3415), .B1(n8023), .C0(n7550), 
        .C1(n8021), .Y(N28078) );
  OAI222XL U12939 ( .A0(n7402), .A1(n8040), .B0(n3347), .B1(n8037), .C0(n7550), 
        .C1(n8034), .Y(N28142) );
  OAI222XL U12940 ( .A0(n7402), .A1(n8077), .B0(n3134), .B1(n8074), .C0(n7550), 
        .C1(n8072), .Y(N28334) );
  OAI222XL U12941 ( .A0(n7402), .A1(n8091), .B0(n3063), .B1(n8087), .C0(n7550), 
        .C1(n8084), .Y(N28398) );
  OAI222XL U12942 ( .A0(n7402), .A1(n8156), .B0(n2580), .B1(n8151), .C0(n7550), 
        .C1(n8148), .Y(N28718) );
  OAI222XL U12943 ( .A0(n7402), .A1(n6588), .B0(n8164), .B1(n2482), .C0(n8162), 
        .C1(n7550), .Y(N28782) );
  OAI222XL U12944 ( .A0(n7404), .A1(n8003), .B0(n3551), .B1(n7999), .C0(n7549), 
        .C1(n7995), .Y(N27951) );
  OAI222XL U12945 ( .A0(n7404), .A1(n8013), .B0(n3483), .B1(n8012), .C0(n7549), 
        .C1(n8007), .Y(N28015) );
  OAI222XL U12946 ( .A0(n7404), .A1(n8027), .B0(n3414), .B1(n8025), .C0(n7549), 
        .C1(n8021), .Y(N28079) );
  OAI222XL U12947 ( .A0(n7404), .A1(n8040), .B0(n3346), .B1(n8037), .C0(n7549), 
        .C1(n8034), .Y(N28143) );
  OAI222XL U12948 ( .A0(n7404), .A1(n8077), .B0(n3133), .B1(n8074), .C0(n7549), 
        .C1(n8072), .Y(N28335) );
  OAI222XL U12949 ( .A0(n7404), .A1(n8091), .B0(n3062), .B1(n8087), .C0(n7549), 
        .C1(n8084), .Y(N28399) );
  OAI222XL U12950 ( .A0(n7404), .A1(n8156), .B0(n2579), .B1(n8152), .C0(n7549), 
        .C1(n8148), .Y(N28719) );
  OAI222XL U12951 ( .A0(n7404), .A1(n6588), .B0(n8165), .B1(n2479), .C0(n8161), 
        .C1(n7549), .Y(N28783) );
  AOI221XL U12952 ( .A0(n8704), .A1(n8157), .B0(n8705), .B1(n8144), .C0(n4617), 
        .Y(n4605) );
  CLKINVX1 U12953 ( .A(n2485), .Y(n8704) );
  CLKINVX1 U12954 ( .A(n2581), .Y(n8705) );
  OAI222XL U12955 ( .A0(n8080), .A1(n3064), .B0(n8016), .B1(n3416), .C0(n8068), 
        .C1(n3135), .Y(n4617) );
  AOI221XL U12956 ( .A0(n8699), .A1(n8157), .B0(n8700), .B1(n8144), .C0(n4599), 
        .Y(n4587) );
  CLKINVX1 U12957 ( .A(n2482), .Y(n8699) );
  CLKINVX1 U12958 ( .A(n2580), .Y(n8700) );
  OAI222XL U12959 ( .A0(n8081), .A1(n3063), .B0(n8017), .B1(n3415), .C0(n8067), 
        .C1(n3134), .Y(n4599) );
  AOI221XL U12960 ( .A0(n8694), .A1(n8157), .B0(n8695), .B1(n8145), .C0(n4581), 
        .Y(n4569) );
  CLKINVX1 U12961 ( .A(n2479), .Y(n8694) );
  CLKINVX1 U12962 ( .A(n2579), .Y(n8695) );
  OAI222XL U12963 ( .A0(n8081), .A1(n3062), .B0(n8017), .B1(n3414), .C0(n8067), 
        .C1(n3133), .Y(n4581) );
  CLKINVX1 U12964 ( .A(n3552), .Y(n8701) );
  CLKINVX1 U12965 ( .A(n3347), .Y(n8702) );
  OAI222XL U12966 ( .A0(n8698), .A1(n7932), .B0(n7929), .B1(n9288), .C0(n8005), 
        .C1(n3484), .Y(n4596) );
  CLKINVX1 U12967 ( .A(n3551), .Y(n8696) );
  CLKINVX1 U12968 ( .A(n3346), .Y(n8697) );
  OAI222XL U12969 ( .A0(n8693), .A1(n7932), .B0(n3676), .B1(n9280), .C0(n8005), 
        .C1(n3483), .Y(n4578) );
  CLKINVX1 U12970 ( .A(n3550), .Y(n8691) );
  CLKINVX1 U12971 ( .A(n3345), .Y(n8692) );
  OAI222XL U12972 ( .A0(n8688), .A1(n3675), .B0(n7931), .B1(n9272), .C0(n8005), 
        .C1(n3482), .Y(n4560) );
  OAI221XL U12973 ( .A0(n7400), .A1(n6584), .B0(n7551), .B1(n7985), .C0(n3623), 
        .Y(N27885) );
  OAI221XL U12974 ( .A0(n7400), .A1(n6583), .B0(n7551), .B1(n8049), .C0(n3277), 
        .Y(N28205) );
  OAI221XL U12975 ( .A0(n7400), .A1(n6605), .B0(n7551), .B1(n8100), .C0(n2994), 
        .Y(N28461) );
  OAI221XL U12976 ( .A0(n7400), .A1(n6606), .B0(n7551), .B1(n8113), .C0(n2909), 
        .Y(N28525) );
  OAI221XL U12977 ( .A0(n7400), .A1(n8130), .B0(n7551), .B1(n8126), .C0(n2787), 
        .Y(N28589) );
  OAI221XL U12978 ( .A0(n7400), .A1(n7976), .B0(n7551), .B1(n7972), .C0(n4603), 
        .Y(N27821) );
  OAI221XL U12979 ( .A0(n7402), .A1(n7988), .B0(n7550), .B1(n7985), .C0(n3622), 
        .Y(N27886) );
  OAI221XL U12980 ( .A0(n7402), .A1(n6583), .B0(n7550), .B1(n8049), .C0(n3276), 
        .Y(N28206) );
  OAI221XL U12981 ( .A0(n7402), .A1(n6605), .B0(n7550), .B1(n8100), .C0(n2993), 
        .Y(N28462) );
  OAI221XL U12982 ( .A0(n7402), .A1(n6606), .B0(n7550), .B1(n8113), .C0(n2907), 
        .Y(N28526) );
  OAI221XL U12983 ( .A0(n7402), .A1(n8130), .B0(n7550), .B1(n8126), .C0(n2786), 
        .Y(N28590) );
  OAI221XL U12984 ( .A0(n7402), .A1(n7976), .B0(n7550), .B1(n7972), .C0(n4585), 
        .Y(N27822) );
  OAI221XL U12985 ( .A0(n7404), .A1(n7988), .B0(n7549), .B1(n7985), .C0(n3621), 
        .Y(N27887) );
  OAI221XL U12986 ( .A0(n7404), .A1(n8052), .B0(n7549), .B1(n8049), .C0(n3275), 
        .Y(N28207) );
  OAI221XL U12987 ( .A0(n7404), .A1(n6605), .B0(n7549), .B1(n8100), .C0(n2992), 
        .Y(N28463) );
  OAI221XL U12988 ( .A0(n7404), .A1(n8116), .B0(n7549), .B1(n8113), .C0(n2905), 
        .Y(N28527) );
  OAI221XL U12989 ( .A0(n7404), .A1(n8130), .B0(n7549), .B1(n8126), .C0(n2785), 
        .Y(N28591) );
  OAI221XL U12990 ( .A0(n7404), .A1(n7976), .B0(n7549), .B1(n7972), .C0(n4567), 
        .Y(N27823) );
  OAI221XL U12991 ( .A0(n7406), .A1(n7988), .B0(n7548), .B1(n7985), .C0(n3620), 
        .Y(N27888) );
  OAI221XL U12992 ( .A0(n7406), .A1(n8052), .B0(n7548), .B1(n8049), .C0(n3274), 
        .Y(N28208) );
  OAI221XL U12993 ( .A0(n7406), .A1(n8103), .B0(n7548), .B1(n8100), .C0(n2991), 
        .Y(N28464) );
  OAI221XL U12994 ( .A0(n7406), .A1(n8116), .B0(n7548), .B1(n8113), .C0(n2903), 
        .Y(N28528) );
  OAI221XL U12995 ( .A0(n7406), .A1(n8130), .B0(n7548), .B1(n8126), .C0(n2784), 
        .Y(N28592) );
  OAI221XL U12996 ( .A0(n7406), .A1(n7976), .B0(n7548), .B1(n7972), .C0(n4549), 
        .Y(N27824) );
  CLKINVX1 U12997 ( .A(n3348), .Y(n8707) );
  CLKINVX1 U12998 ( .A(n3553), .Y(n8706) );
  CLKBUFX3 U12999 ( .A(n8411), .Y(n7006) );
  CLKBUFX3 U13000 ( .A(n8412), .Y(n7004) );
  CLKBUFX3 U13001 ( .A(n7001), .Y(n6991) );
  CLKBUFX3 U13002 ( .A(n8413), .Y(n7001) );
  OAI222XL U13003 ( .A0(n9322), .A1(n7943), .B0(n8718), .B1(n7938), .C0(n7935), 
        .C1(n9321), .Y(n4665) );
  OAI222XL U13004 ( .A0(n7957), .A1(n9319), .B0(n9326), .B1(n7954), .C0(n8718), 
        .C1(n7951), .Y(n4663) );
  OAI222XL U13005 ( .A0(n9314), .A1(n7943), .B0(n8713), .B1(n7939), .C0(n7935), 
        .C1(n9313), .Y(n4647) );
  OAI222XL U13006 ( .A0(n7958), .A1(n9311), .B0(n9318), .B1(n7954), .C0(n8713), 
        .C1(n7951), .Y(n4645) );
  OAI222XL U13007 ( .A0(n8708), .A1(n7933), .B0(n7929), .B1(n9304), .C0(n8004), 
        .C1(n3486), .Y(n4632) );
  OAI222XL U13008 ( .A0(n7956), .A1(n9303), .B0(n9310), .B1(n7954), .C0(n8708), 
        .C1(n7951), .Y(n4627) );
  OAI222XL U13009 ( .A0(n7392), .A1(n8001), .B0(n3557), .B1(n7998), .C0(n7555), 
        .C1(n7996), .Y(N27945) );
  OAI222XL U13010 ( .A0(n7392), .A1(n8015), .B0(n3489), .B1(n8011), .C0(n7555), 
        .C1(n6618), .Y(N28009) );
  OAI222XL U13011 ( .A0(n7392), .A1(n8026), .B0(n3420), .B1(n8024), .C0(n7555), 
        .C1(n8020), .Y(N28073) );
  OAI222XL U13012 ( .A0(n7392), .A1(n8039), .B0(n3352), .B1(n8038), .C0(n7555), 
        .C1(n8033), .Y(N28137) );
  OAI222XL U13013 ( .A0(n7392), .A1(n8078), .B0(n3139), .B1(n8076), .C0(n7555), 
        .C1(n8071), .Y(N28329) );
  OAI222XL U13014 ( .A0(n7392), .A1(n8090), .B0(n3068), .B1(n8088), .C0(n7555), 
        .C1(n8086), .Y(N28393) );
  OAI222XL U13015 ( .A0(n7392), .A1(n8154), .B0(n2585), .B1(n8152), .C0(n7555), 
        .C1(n6615), .Y(N28713) );
  OAI222XL U13016 ( .A0(n7392), .A1(n8169), .B0(n8166), .B1(n2497), .C0(n8162), 
        .C1(n7555), .Y(N28777) );
  OAI222XL U13017 ( .A0(n7394), .A1(n8001), .B0(n3556), .B1(n7998), .C0(n7554), 
        .C1(n6617), .Y(N27946) );
  OAI222XL U13018 ( .A0(n7394), .A1(n3431), .B0(n3488), .B1(n6589), .C0(n7554), 
        .C1(n6618), .Y(N28010) );
  OAI222XL U13019 ( .A0(n7394), .A1(n8026), .B0(n3419), .B1(n8023), .C0(n7554), 
        .C1(n8020), .Y(N28074) );
  OAI222XL U13020 ( .A0(n7394), .A1(n8039), .B0(n3351), .B1(n8036), .C0(n7554), 
        .C1(n8033), .Y(N28138) );
  OAI222XL U13021 ( .A0(n7394), .A1(n3081), .B0(n3138), .B1(n6590), .C0(n7554), 
        .C1(n8071), .Y(N28330) );
  OAI222XL U13022 ( .A0(n7394), .A1(n8090), .B0(n3067), .B1(n8089), .C0(n7554), 
        .C1(n6619), .Y(N28394) );
  OAI222XL U13023 ( .A0(n7394), .A1(n8154), .B0(n2584), .B1(n8153), .C0(n7554), 
        .C1(n6615), .Y(N28714) );
  OAI222XL U13024 ( .A0(n7394), .A1(n8169), .B0(n8166), .B1(n2494), .C0(n8162), 
        .C1(n7554), .Y(N28778) );
  OAI222XL U13025 ( .A0(n7396), .A1(n8001), .B0(n3555), .B1(n8000), .C0(n7553), 
        .C1(n6617), .Y(N27947) );
  OAI222XL U13026 ( .A0(n7396), .A1(n3431), .B0(n3487), .B1(n6589), .C0(n7553), 
        .C1(n6618), .Y(N28011) );
  OAI222XL U13027 ( .A0(n7396), .A1(n8026), .B0(n3418), .B1(n6577), .C0(n7553), 
        .C1(n8020), .Y(N28075) );
  OAI222XL U13028 ( .A0(n7396), .A1(n8039), .B0(n3350), .B1(n8036), .C0(n7553), 
        .C1(n8033), .Y(N28139) );
  OAI222XL U13029 ( .A0(n7396), .A1(n3081), .B0(n3137), .B1(n6590), .C0(n7553), 
        .C1(n8071), .Y(N28331) );
  OAI222XL U13030 ( .A0(n7396), .A1(n8090), .B0(n3066), .B1(n8089), .C0(n7553), 
        .C1(n6619), .Y(N28395) );
  OAI222XL U13031 ( .A0(n7396), .A1(n8154), .B0(n2583), .B1(n8153), .C0(n7553), 
        .C1(n6615), .Y(N28715) );
  OAI222XL U13032 ( .A0(n7396), .A1(n8169), .B0(n8166), .B1(n2491), .C0(n8162), 
        .C1(n7553), .Y(N28779) );
  OAI222XL U13033 ( .A0(n7398), .A1(n8001), .B0(n3554), .B1(n7999), .C0(n7552), 
        .C1(n6617), .Y(N27948) );
  OAI222XL U13034 ( .A0(n7398), .A1(n3431), .B0(n3486), .B1(n6589), .C0(n7552), 
        .C1(n6618), .Y(N28012) );
  OAI222XL U13035 ( .A0(n7398), .A1(n8026), .B0(n3417), .B1(n6577), .C0(n7552), 
        .C1(n8020), .Y(N28076) );
  OAI222XL U13036 ( .A0(n7398), .A1(n8039), .B0(n3349), .B1(n6575), .C0(n7552), 
        .C1(n8033), .Y(N28140) );
  OAI222XL U13037 ( .A0(n7398), .A1(n3081), .B0(n3136), .B1(n6590), .C0(n7552), 
        .C1(n8071), .Y(N28332) );
  OAI222XL U13038 ( .A0(n7398), .A1(n8090), .B0(n3065), .B1(n6578), .C0(n7552), 
        .C1(n6619), .Y(N28396) );
  OAI222XL U13039 ( .A0(n7398), .A1(n8154), .B0(n2582), .B1(n8151), .C0(n7552), 
        .C1(n6615), .Y(N28716) );
  OAI222XL U13040 ( .A0(n7398), .A1(n8169), .B0(n8166), .B1(n2488), .C0(n8162), 
        .C1(n7552), .Y(N28780) );
  AOI221XL U13041 ( .A0(n8724), .A1(n8160), .B0(n8725), .B1(n8144), .C0(n4689), 
        .Y(n4677) );
  CLKINVX1 U13042 ( .A(n2497), .Y(n8724) );
  CLKINVX1 U13043 ( .A(n2585), .Y(n8725) );
  OAI222XL U13044 ( .A0(n8080), .A1(n3068), .B0(n8016), .B1(n3420), .C0(n8068), 
        .C1(n3139), .Y(n4689) );
  AOI221XL U13045 ( .A0(n8719), .A1(n8157), .B0(n8720), .B1(n8144), .C0(n4671), 
        .Y(n4659) );
  CLKINVX1 U13046 ( .A(n2494), .Y(n8719) );
  CLKINVX1 U13047 ( .A(n2584), .Y(n8720) );
  OAI222XL U13048 ( .A0(n8080), .A1(n3067), .B0(n8016), .B1(n3419), .C0(n8068), 
        .C1(n3138), .Y(n4671) );
  AOI221XL U13049 ( .A0(n8714), .A1(n8157), .B0(n8715), .B1(n8144), .C0(n4653), 
        .Y(n4641) );
  CLKINVX1 U13050 ( .A(n2491), .Y(n8714) );
  CLKINVX1 U13051 ( .A(n2583), .Y(n8715) );
  OAI222XL U13052 ( .A0(n8080), .A1(n3066), .B0(n8016), .B1(n3418), .C0(n8068), 
        .C1(n3137), .Y(n4653) );
  AOI221XL U13053 ( .A0(n8709), .A1(n8157), .B0(n8710), .B1(n8144), .C0(n4635), 
        .Y(n4623) );
  CLKINVX1 U13054 ( .A(n2488), .Y(n8709) );
  CLKINVX1 U13055 ( .A(n2582), .Y(n8710) );
  OAI222XL U13056 ( .A0(n8080), .A1(n3065), .B0(n8016), .B1(n3417), .C0(n8068), 
        .C1(n3136), .Y(n4635) );
  CLKINVX1 U13057 ( .A(n3557), .Y(n8726) );
  CLKINVX1 U13058 ( .A(n3352), .Y(n8727) );
  OAI222XL U13059 ( .A0(n8723), .A1(n7932), .B0(n7929), .B1(n9328), .C0(n8004), 
        .C1(n3489), .Y(n4686) );
  CLKINVX1 U13060 ( .A(n3556), .Y(n8721) );
  CLKINVX1 U13061 ( .A(n3351), .Y(n8722) );
  OAI222XL U13062 ( .A0(n8718), .A1(n7932), .B0(n7929), .B1(n9320), .C0(n8004), 
        .C1(n3488), .Y(n4668) );
  CLKINVX1 U13063 ( .A(n3555), .Y(n8716) );
  CLKINVX1 U13064 ( .A(n3350), .Y(n8717) );
  OAI222XL U13065 ( .A0(n8713), .A1(n7932), .B0(n7929), .B1(n9312), .C0(n8004), 
        .C1(n3487), .Y(n4650) );
  OAI221XL U13066 ( .A0(n7392), .A1(n7989), .B0(n7555), .B1(n7986), .C0(n3627), 
        .Y(N27881) );
  OAI221XL U13067 ( .A0(n7392), .A1(n8053), .B0(n7555), .B1(n8050), .C0(n3281), 
        .Y(N28201) );
  OAI221XL U13068 ( .A0(n7392), .A1(n8104), .B0(n7555), .B1(n8101), .C0(n2998), 
        .Y(N28457) );
  OAI221XL U13069 ( .A0(n7392), .A1(n8117), .B0(n7555), .B1(n8114), .C0(n2917), 
        .Y(N28521) );
  OAI221XL U13070 ( .A0(n7392), .A1(n8129), .B0(n7555), .B1(n8127), .C0(n2791), 
        .Y(N28585) );
  OAI221XL U13071 ( .A0(n7392), .A1(n7975), .B0(n7555), .B1(n7973), .C0(n4675), 
        .Y(N27817) );
  OAI221XL U13072 ( .A0(n7394), .A1(n7989), .B0(n7554), .B1(n7986), .C0(n3626), 
        .Y(N27882) );
  OAI221XL U13073 ( .A0(n7394), .A1(n8053), .B0(n7554), .B1(n8050), .C0(n3280), 
        .Y(N28202) );
  OAI221XL U13074 ( .A0(n7394), .A1(n8104), .B0(n7554), .B1(n8101), .C0(n2997), 
        .Y(N28458) );
  OAI221XL U13075 ( .A0(n7394), .A1(n8117), .B0(n7554), .B1(n8114), .C0(n2915), 
        .Y(N28522) );
  OAI221XL U13076 ( .A0(n7394), .A1(n8129), .B0(n7554), .B1(n8127), .C0(n2790), 
        .Y(N28586) );
  OAI221XL U13077 ( .A0(n7394), .A1(n7975), .B0(n7554), .B1(n7973), .C0(n4657), 
        .Y(N27818) );
  OAI221XL U13078 ( .A0(n7396), .A1(n7989), .B0(n7553), .B1(n7986), .C0(n3625), 
        .Y(N27883) );
  OAI221XL U13079 ( .A0(n7396), .A1(n8053), .B0(n7553), .B1(n8050), .C0(n3279), 
        .Y(N28203) );
  OAI221XL U13080 ( .A0(n7396), .A1(n8104), .B0(n7553), .B1(n8101), .C0(n2996), 
        .Y(N28459) );
  OAI221XL U13081 ( .A0(n7396), .A1(n8117), .B0(n7553), .B1(n8114), .C0(n2913), 
        .Y(N28523) );
  OAI221XL U13082 ( .A0(n7396), .A1(n8129), .B0(n7553), .B1(n8127), .C0(n2789), 
        .Y(N28587) );
  OAI221XL U13083 ( .A0(n7396), .A1(n7975), .B0(n7553), .B1(n7973), .C0(n4639), 
        .Y(N27819) );
  OAI221XL U13084 ( .A0(n7398), .A1(n7989), .B0(n7552), .B1(n7986), .C0(n3624), 
        .Y(N27884) );
  OAI221XL U13085 ( .A0(n7398), .A1(n8053), .B0(n7552), .B1(n8050), .C0(n3278), 
        .Y(N28204) );
  OAI221XL U13086 ( .A0(n7398), .A1(n8104), .B0(n7552), .B1(n8101), .C0(n2995), 
        .Y(N28460) );
  OAI221XL U13087 ( .A0(n7398), .A1(n8117), .B0(n7552), .B1(n8114), .C0(n2911), 
        .Y(N28524) );
  OAI221XL U13088 ( .A0(n7398), .A1(n8129), .B0(n7552), .B1(n8127), .C0(n2788), 
        .Y(N28588) );
  OAI221XL U13089 ( .A0(n7398), .A1(n7975), .B0(n7552), .B1(n7973), .C0(n4621), 
        .Y(N27820) );
  CLKINVX1 U13090 ( .A(n3349), .Y(n8712) );
  CLKINVX1 U13091 ( .A(n3554), .Y(n8711) );
  OAI222XL U13092 ( .A0(n9370), .A1(n3669), .B0(n8748), .B1(n7938), .C0(n7935), 
        .C1(n9369), .Y(n4773) );
  OAI222XL U13093 ( .A0(n7956), .A1(n9367), .B0(n9374), .B1(n7955), .C0(n8748), 
        .C1(n7950), .Y(n4771) );
  OAI222XL U13094 ( .A0(n9362), .A1(n7943), .B0(n8743), .B1(n7940), .C0(n7935), 
        .C1(n9361), .Y(n4755) );
  OAI222XL U13095 ( .A0(n7956), .A1(n9359), .B0(n9366), .B1(n7954), .C0(n8743), 
        .C1(n3665), .Y(n4753) );
  OAI222XL U13096 ( .A0(n9354), .A1(n7943), .B0(n8738), .B1(n7939), .C0(n7935), 
        .C1(n9353), .Y(n4737) );
  OAI222XL U13097 ( .A0(n7956), .A1(n9351), .B0(n9358), .B1(n7954), .C0(n8738), 
        .C1(n7951), .Y(n4735) );
  OAI222XL U13098 ( .A0(n9346), .A1(n7943), .B0(n8733), .B1(n7938), .C0(n7935), 
        .C1(n9345), .Y(n4719) );
  OAI222XL U13099 ( .A0(n7958), .A1(n9343), .B0(n9350), .B1(n7954), .C0(n8733), 
        .C1(n7951), .Y(n4717) );
  OAI222XL U13100 ( .A0(n9338), .A1(n7943), .B0(n8728), .B1(n7939), .C0(n7935), 
        .C1(n9337), .Y(n4701) );
  OAI222XL U13101 ( .A0(n7956), .A1(n9335), .B0(n9342), .B1(n7954), .C0(n8728), 
        .C1(n7950), .Y(n4699) );
  OAI222XL U13102 ( .A0(n9330), .A1(n7943), .B0(n8723), .B1(n7938), .C0(n7935), 
        .C1(n9329), .Y(n4683) );
  OAI222XL U13103 ( .A0(n7957), .A1(n9327), .B0(n9334), .B1(n7954), .C0(n8723), 
        .C1(n7952), .Y(n4681) );
  OAI222XL U13104 ( .A0(n7380), .A1(n8001), .B0(n3563), .B1(n8000), .C0(n7561), 
        .C1(n7997), .Y(N27939) );
  OAI222XL U13105 ( .A0(n7380), .A1(n3431), .B0(n3495), .B1(n8010), .C0(n7561), 
        .C1(n8008), .Y(N28003) );
  OAI222XL U13106 ( .A0(n7380), .A1(n8026), .B0(n3426), .B1(n6577), .C0(n7561), 
        .C1(n8020), .Y(N28067) );
  OAI222XL U13107 ( .A0(n7380), .A1(n8039), .B0(n3358), .B1(n8038), .C0(n7561), 
        .C1(n8033), .Y(N28131) );
  OAI222XL U13108 ( .A0(n7380), .A1(n8078), .B0(n3145), .B1(n8074), .C0(n7561), 
        .C1(n8071), .Y(N28323) );
  OAI222XL U13109 ( .A0(n7380), .A1(n8090), .B0(n3074), .B1(n6578), .C0(n7561), 
        .C1(n6619), .Y(N28387) );
  OAI222XL U13110 ( .A0(n7380), .A1(n8154), .B0(n2591), .B1(n8153), .C0(n7561), 
        .C1(n8149), .Y(N28707) );
  OAI222XL U13111 ( .A0(n7380), .A1(n8169), .B0(n8166), .B1(n2515), .C0(n8162), 
        .C1(n7561), .Y(N28771) );
  OAI222XL U13112 ( .A0(n7382), .A1(n8001), .B0(n3562), .B1(n8000), .C0(n7560), 
        .C1(n7996), .Y(N27940) );
  OAI222XL U13113 ( .A0(n7382), .A1(n8014), .B0(n3494), .B1(n8011), .C0(n7560), 
        .C1(n8009), .Y(N28004) );
  OAI222XL U13114 ( .A0(n7382), .A1(n8026), .B0(n3425), .B1(n8024), .C0(n7560), 
        .C1(n8020), .Y(N28068) );
  OAI222XL U13115 ( .A0(n7382), .A1(n8039), .B0(n3357), .B1(n6575), .C0(n7560), 
        .C1(n8033), .Y(N28132) );
  OAI222XL U13116 ( .A0(n7382), .A1(n8079), .B0(n3144), .B1(n8076), .C0(n7560), 
        .C1(n8071), .Y(N28324) );
  OAI222XL U13117 ( .A0(n7382), .A1(n8090), .B0(n3073), .B1(n8088), .C0(n7560), 
        .C1(n8085), .Y(N28388) );
  OAI222XL U13118 ( .A0(n7382), .A1(n8154), .B0(n2590), .B1(n8152), .C0(n7560), 
        .C1(n8150), .Y(N28708) );
  OAI222XL U13119 ( .A0(n7382), .A1(n8169), .B0(n8164), .B1(n2512), .C0(n8162), 
        .C1(n7560), .Y(N28772) );
  OAI222XL U13120 ( .A0(n7384), .A1(n8001), .B0(n3561), .B1(n6581), .C0(n7559), 
        .C1(n7997), .Y(N27941) );
  OAI222XL U13121 ( .A0(n7384), .A1(n8014), .B0(n3493), .B1(n8011), .C0(n7559), 
        .C1(n8008), .Y(N28005) );
  OAI222XL U13122 ( .A0(n7384), .A1(n8026), .B0(n3424), .B1(n8024), .C0(n7559), 
        .C1(n8020), .Y(N28069) );
  OAI222XL U13123 ( .A0(n7384), .A1(n8039), .B0(n3356), .B1(n8038), .C0(n7559), 
        .C1(n8033), .Y(N28133) );
  OAI222XL U13124 ( .A0(n7384), .A1(n8079), .B0(n3143), .B1(n8076), .C0(n7559), 
        .C1(n8071), .Y(N28325) );
  OAI222XL U13125 ( .A0(n7384), .A1(n8090), .B0(n3072), .B1(n8088), .C0(n7559), 
        .C1(n8086), .Y(N28389) );
  OAI222XL U13126 ( .A0(n7384), .A1(n8154), .B0(n2589), .B1(n6587), .C0(n7559), 
        .C1(n8149), .Y(N28709) );
  OAI222XL U13127 ( .A0(n7384), .A1(n8169), .B0(n8164), .B1(n2509), .C0(n8162), 
        .C1(n7559), .Y(N28773) );
  OAI222XL U13128 ( .A0(n7386), .A1(n8001), .B0(n3560), .B1(n8000), .C0(n7558), 
        .C1(n7996), .Y(N27942) );
  OAI222XL U13129 ( .A0(n7386), .A1(n8015), .B0(n3492), .B1(n8011), .C0(n7558), 
        .C1(n8009), .Y(N28006) );
  OAI222XL U13130 ( .A0(n7386), .A1(n8026), .B0(n3423), .B1(n8024), .C0(n7558), 
        .C1(n8020), .Y(N28070) );
  OAI222XL U13131 ( .A0(n7386), .A1(n8039), .B0(n3355), .B1(n8037), .C0(n7558), 
        .C1(n8033), .Y(N28134) );
  OAI222XL U13132 ( .A0(n7386), .A1(n8078), .B0(n3142), .B1(n8075), .C0(n7558), 
        .C1(n8071), .Y(N28326) );
  OAI222XL U13133 ( .A0(n7386), .A1(n8090), .B0(n3071), .B1(n8087), .C0(n7558), 
        .C1(n8085), .Y(N28390) );
  OAI222XL U13134 ( .A0(n7386), .A1(n8154), .B0(n2588), .B1(n8153), .C0(n7558), 
        .C1(n8150), .Y(N28710) );
  OAI222XL U13135 ( .A0(n7386), .A1(n8169), .B0(n8164), .B1(n2506), .C0(n8162), 
        .C1(n7558), .Y(N28774) );
  OAI222XL U13136 ( .A0(n7388), .A1(n8001), .B0(n3559), .B1(n7999), .C0(n7557), 
        .C1(n7997), .Y(N27943) );
  OAI222XL U13137 ( .A0(n7388), .A1(n8014), .B0(n3491), .B1(n8012), .C0(n7557), 
        .C1(n8008), .Y(N28007) );
  OAI222XL U13138 ( .A0(n7388), .A1(n8026), .B0(n3422), .B1(n8023), .C0(n7557), 
        .C1(n8020), .Y(N28071) );
  OAI222XL U13139 ( .A0(n7388), .A1(n8039), .B0(n3354), .B1(n8036), .C0(n7557), 
        .C1(n8033), .Y(N28135) );
  OAI222XL U13140 ( .A0(n7388), .A1(n8079), .B0(n3141), .B1(n8074), .C0(n7557), 
        .C1(n8071), .Y(N28327) );
  OAI222XL U13141 ( .A0(n7388), .A1(n8090), .B0(n3070), .B1(n8089), .C0(n7557), 
        .C1(n8086), .Y(N28391) );
  OAI222XL U13142 ( .A0(n7388), .A1(n8154), .B0(n2587), .B1(n8151), .C0(n7557), 
        .C1(n8149), .Y(N28711) );
  OAI222XL U13143 ( .A0(n7388), .A1(n8169), .B0(n8166), .B1(n2503), .C0(n8162), 
        .C1(n7557), .Y(N28775) );
  OAI222XL U13144 ( .A0(n7390), .A1(n8001), .B0(n3558), .B1(n7998), .C0(n7556), 
        .C1(n7996), .Y(N27944) );
  OAI222XL U13145 ( .A0(n7390), .A1(n8015), .B0(n3490), .B1(n8010), .C0(n7556), 
        .C1(n8009), .Y(N28008) );
  OAI222XL U13146 ( .A0(n7390), .A1(n8026), .B0(n3421), .B1(n8025), .C0(n7556), 
        .C1(n8020), .Y(N28072) );
  OAI222XL U13147 ( .A0(n7390), .A1(n8039), .B0(n3353), .B1(n8038), .C0(n7556), 
        .C1(n8033), .Y(N28136) );
  OAI222XL U13148 ( .A0(n7390), .A1(n3081), .B0(n3140), .B1(n8076), .C0(n7556), 
        .C1(n8071), .Y(N28328) );
  OAI222XL U13149 ( .A0(n7390), .A1(n8090), .B0(n3069), .B1(n8088), .C0(n7556), 
        .C1(n8085), .Y(N28392) );
  OAI222XL U13150 ( .A0(n7390), .A1(n8154), .B0(n2586), .B1(n8152), .C0(n7556), 
        .C1(n8150), .Y(N28712) );
  OAI222XL U13151 ( .A0(n7390), .A1(n8169), .B0(n8166), .B1(n2500), .C0(n8162), 
        .C1(n7556), .Y(N28776) );
  AOI221XL U13152 ( .A0(n8754), .A1(n8159), .B0(n8755), .B1(n8144), .C0(n4797), 
        .Y(n4785) );
  CLKINVX1 U13153 ( .A(n2515), .Y(n8754) );
  CLKINVX1 U13154 ( .A(n2591), .Y(n8755) );
  OAI222XL U13155 ( .A0(n8082), .A1(n3074), .B0(n8016), .B1(n3426), .C0(n8068), 
        .C1(n3145), .Y(n4797) );
  AOI221XL U13156 ( .A0(n8749), .A1(n8157), .B0(n8750), .B1(n8144), .C0(n4779), 
        .Y(n4767) );
  CLKINVX1 U13157 ( .A(n2512), .Y(n8749) );
  CLKINVX1 U13158 ( .A(n2590), .Y(n8750) );
  OAI222XL U13159 ( .A0(n8082), .A1(n3073), .B0(n8016), .B1(n3425), .C0(n8068), 
        .C1(n3144), .Y(n4779) );
  AOI221XL U13160 ( .A0(n8744), .A1(n6610), .B0(n8745), .B1(n8144), .C0(n4761), 
        .Y(n4749) );
  CLKINVX1 U13161 ( .A(n2509), .Y(n8744) );
  CLKINVX1 U13162 ( .A(n2589), .Y(n8745) );
  OAI222XL U13163 ( .A0(n8080), .A1(n3072), .B0(n8016), .B1(n3424), .C0(n8068), 
        .C1(n3143), .Y(n4761) );
  AOI221XL U13164 ( .A0(n8739), .A1(n6610), .B0(n8740), .B1(n8144), .C0(n4743), 
        .Y(n4731) );
  CLKINVX1 U13165 ( .A(n2506), .Y(n8739) );
  CLKINVX1 U13166 ( .A(n2588), .Y(n8740) );
  OAI222XL U13167 ( .A0(n8082), .A1(n3071), .B0(n8016), .B1(n3423), .C0(n8068), 
        .C1(n3142), .Y(n4743) );
  AOI221XL U13168 ( .A0(n8734), .A1(n6610), .B0(n8735), .B1(n8144), .C0(n4725), 
        .Y(n4713) );
  CLKINVX1 U13169 ( .A(n2503), .Y(n8734) );
  CLKINVX1 U13170 ( .A(n2587), .Y(n8735) );
  OAI222XL U13171 ( .A0(n8082), .A1(n3070), .B0(n8016), .B1(n3422), .C0(n8068), 
        .C1(n3141), .Y(n4725) );
  AOI221XL U13172 ( .A0(n8729), .A1(n8159), .B0(n8730), .B1(n8144), .C0(n4707), 
        .Y(n4695) );
  CLKINVX1 U13173 ( .A(n2500), .Y(n8729) );
  CLKINVX1 U13174 ( .A(n2586), .Y(n8730) );
  OAI222XL U13175 ( .A0(n8082), .A1(n3069), .B0(n8016), .B1(n3421), .C0(n8068), 
        .C1(n3140), .Y(n4707) );
  CLKINVX1 U13176 ( .A(n3563), .Y(n8756) );
  CLKINVX1 U13177 ( .A(n3358), .Y(n8757) );
  OAI222XL U13178 ( .A0(n8753), .A1(n7934), .B0(n7929), .B1(n9376), .C0(n8004), 
        .C1(n3495), .Y(n4794) );
  CLKINVX1 U13179 ( .A(n3562), .Y(n8751) );
  CLKINVX1 U13180 ( .A(n3357), .Y(n8752) );
  OAI222XL U13181 ( .A0(n8748), .A1(n7934), .B0(n7929), .B1(n9368), .C0(n8004), 
        .C1(n3494), .Y(n4776) );
  CLKINVX1 U13182 ( .A(n3561), .Y(n8746) );
  CLKINVX1 U13183 ( .A(n3356), .Y(n8747) );
  OAI222XL U13184 ( .A0(n8743), .A1(n7933), .B0(n7931), .B1(n9360), .C0(n8004), 
        .C1(n3493), .Y(n4758) );
  CLKINVX1 U13185 ( .A(n3560), .Y(n8741) );
  CLKINVX1 U13186 ( .A(n3355), .Y(n8742) );
  OAI222XL U13187 ( .A0(n8738), .A1(n7932), .B0(n7929), .B1(n9352), .C0(n8004), 
        .C1(n3492), .Y(n4740) );
  CLKINVX1 U13188 ( .A(n3559), .Y(n8736) );
  CLKINVX1 U13189 ( .A(n3354), .Y(n8737) );
  OAI222XL U13190 ( .A0(n8733), .A1(n7933), .B0(n7929), .B1(n9344), .C0(n8004), 
        .C1(n3491), .Y(n4722) );
  CLKINVX1 U13191 ( .A(n3558), .Y(n8731) );
  CLKINVX1 U13192 ( .A(n3353), .Y(n8732) );
  OAI222XL U13193 ( .A0(n8728), .A1(n7933), .B0(n7929), .B1(n9336), .C0(n8004), 
        .C1(n3490), .Y(n4704) );
  OAI221XL U13194 ( .A0(n7380), .A1(n7989), .B0(n7561), .B1(n7986), .C0(n3633), 
        .Y(N27875) );
  OAI221XL U13195 ( .A0(n7380), .A1(n8053), .B0(n7561), .B1(n8050), .C0(n3287), 
        .Y(N28195) );
  OAI221XL U13196 ( .A0(n7380), .A1(n8104), .B0(n7561), .B1(n8101), .C0(n3004), 
        .Y(N28451) );
  OAI221XL U13197 ( .A0(n7380), .A1(n8117), .B0(n7561), .B1(n8114), .C0(n2929), 
        .Y(N28515) );
  OAI221XL U13198 ( .A0(n7380), .A1(n8129), .B0(n7561), .B1(n8127), .C0(n2797), 
        .Y(N28579) );
  OAI221XL U13199 ( .A0(n7380), .A1(n7975), .B0(n7561), .B1(n7973), .C0(n4783), 
        .Y(N27811) );
  OAI221XL U13200 ( .A0(n7382), .A1(n7989), .B0(n7560), .B1(n7986), .C0(n3632), 
        .Y(N27876) );
  OAI221XL U13201 ( .A0(n7382), .A1(n8053), .B0(n7560), .B1(n8050), .C0(n3286), 
        .Y(N28196) );
  OAI221XL U13202 ( .A0(n7382), .A1(n8104), .B0(n7560), .B1(n8101), .C0(n3003), 
        .Y(N28452) );
  OAI221XL U13203 ( .A0(n7382), .A1(n8117), .B0(n7560), .B1(n8114), .C0(n2927), 
        .Y(N28516) );
  OAI221XL U13204 ( .A0(n7382), .A1(n8129), .B0(n7560), .B1(n8127), .C0(n2796), 
        .Y(N28580) );
  OAI221XL U13205 ( .A0(n7382), .A1(n7975), .B0(n7560), .B1(n7973), .C0(n4765), 
        .Y(N27812) );
  OAI221XL U13206 ( .A0(n7384), .A1(n7989), .B0(n7559), .B1(n7986), .C0(n3631), 
        .Y(N27877) );
  OAI221XL U13207 ( .A0(n7384), .A1(n8053), .B0(n7559), .B1(n8050), .C0(n3285), 
        .Y(N28197) );
  OAI221XL U13208 ( .A0(n7384), .A1(n8104), .B0(n7559), .B1(n8101), .C0(n3002), 
        .Y(N28453) );
  OAI221XL U13209 ( .A0(n7384), .A1(n8117), .B0(n7559), .B1(n8114), .C0(n2925), 
        .Y(N28517) );
  OAI221XL U13210 ( .A0(n7384), .A1(n8129), .B0(n7559), .B1(n8127), .C0(n2795), 
        .Y(N28581) );
  OAI221XL U13211 ( .A0(n7384), .A1(n7975), .B0(n7559), .B1(n7973), .C0(n4747), 
        .Y(N27813) );
  OAI221XL U13212 ( .A0(n7386), .A1(n7989), .B0(n7558), .B1(n7986), .C0(n3630), 
        .Y(N27878) );
  OAI221XL U13213 ( .A0(n7386), .A1(n8053), .B0(n7558), .B1(n8050), .C0(n3284), 
        .Y(N28198) );
  OAI221XL U13214 ( .A0(n7386), .A1(n8104), .B0(n7558), .B1(n8101), .C0(n3001), 
        .Y(N28454) );
  OAI221XL U13215 ( .A0(n7386), .A1(n8117), .B0(n7558), .B1(n8114), .C0(n2923), 
        .Y(N28518) );
  OAI221XL U13216 ( .A0(n7386), .A1(n8129), .B0(n7558), .B1(n8127), .C0(n2794), 
        .Y(N28582) );
  OAI221XL U13217 ( .A0(n7386), .A1(n7975), .B0(n7558), .B1(n7973), .C0(n4729), 
        .Y(N27814) );
  OAI221XL U13218 ( .A0(n7388), .A1(n7989), .B0(n7557), .B1(n7986), .C0(n3629), 
        .Y(N27879) );
  OAI221XL U13219 ( .A0(n7388), .A1(n8053), .B0(n7557), .B1(n8050), .C0(n3283), 
        .Y(N28199) );
  OAI221XL U13220 ( .A0(n7388), .A1(n8104), .B0(n7557), .B1(n8101), .C0(n3000), 
        .Y(N28455) );
  OAI221XL U13221 ( .A0(n7388), .A1(n8117), .B0(n7557), .B1(n8114), .C0(n2921), 
        .Y(N28519) );
  OAI221XL U13222 ( .A0(n7388), .A1(n8129), .B0(n7557), .B1(n8127), .C0(n2793), 
        .Y(N28583) );
  OAI221XL U13223 ( .A0(n7388), .A1(n7975), .B0(n7557), .B1(n7973), .C0(n4711), 
        .Y(N27815) );
  OAI221XL U13224 ( .A0(n7390), .A1(n7989), .B0(n7556), .B1(n7986), .C0(n3628), 
        .Y(N27880) );
  OAI221XL U13225 ( .A0(n7390), .A1(n8053), .B0(n7556), .B1(n8050), .C0(n3282), 
        .Y(N28200) );
  OAI221XL U13226 ( .A0(n7390), .A1(n8104), .B0(n7556), .B1(n8101), .C0(n2999), 
        .Y(N28456) );
  OAI221XL U13227 ( .A0(n7390), .A1(n8117), .B0(n7556), .B1(n8114), .C0(n2919), 
        .Y(N28520) );
  OAI221XL U13228 ( .A0(n7390), .A1(n8129), .B0(n7556), .B1(n8127), .C0(n2792), 
        .Y(N28584) );
  OAI221XL U13229 ( .A0(n7390), .A1(n7975), .B0(n7556), .B1(n7973), .C0(n4693), 
        .Y(N27816) );
  OAI222XL U13230 ( .A0(n8763), .A1(n7934), .B0(n7931), .B1(n9392), .C0(n8006), 
        .C1(n3497), .Y(n4857) );
  OAI222XL U13231 ( .A0(n7956), .A1(n9391), .B0(n9398), .B1(n7955), .C0(n8763), 
        .C1(n7952), .Y(n4838) );
  OAI222XL U13232 ( .A0(n8758), .A1(n7934), .B0(n7929), .B1(n9384), .C0(n8004), 
        .C1(n3496), .Y(n4812) );
  OAI222XL U13233 ( .A0(n7957), .A1(n9383), .B0(n9390), .B1(n7955), .C0(n8758), 
        .C1(n7950), .Y(n4807) );
  OAI222XL U13234 ( .A0(n9378), .A1(n7943), .B0(n8753), .B1(n7939), .C0(n7935), 
        .C1(n9377), .Y(n4791) );
  OAI222XL U13235 ( .A0(n7956), .A1(n9375), .B0(n9382), .B1(n7955), .C0(n8753), 
        .C1(n7950), .Y(n4789) );
  OAI222XL U13236 ( .A0(n7376), .A1(n8001), .B0(n3565), .B1(n6581), .C0(n7563), 
        .C1(n7997), .Y(N27937) );
  OAI222XL U13237 ( .A0(n7376), .A1(n8015), .B0(n3497), .B1(n8011), .C0(n7563), 
        .C1(n8008), .Y(N28001) );
  OAI222XL U13238 ( .A0(n7376), .A1(n8026), .B0(n3428), .B1(n8023), .C0(n7563), 
        .C1(n8020), .Y(N28065) );
  OAI222XL U13239 ( .A0(n7376), .A1(n8039), .B0(n3360), .B1(n8038), .C0(n7563), 
        .C1(n8033), .Y(N28129) );
  OAI222XL U13240 ( .A0(n7376), .A1(n8078), .B0(n3147), .B1(n8075), .C0(n7563), 
        .C1(n8071), .Y(N28321) );
  OAI222XL U13241 ( .A0(n7376), .A1(n8090), .B0(n3076), .B1(n8088), .C0(n7563), 
        .C1(n8085), .Y(N28385) );
  OAI222XL U13242 ( .A0(n7376), .A1(n8154), .B0(n2593), .B1(n8151), .C0(n7563), 
        .C1(n8149), .Y(N28705) );
  OAI222XL U13243 ( .A0(n7376), .A1(n8169), .B0(n8164), .B1(n2521), .C0(n8162), 
        .C1(n7563), .Y(N28769) );
  OAI222XL U13244 ( .A0(n7378), .A1(n8001), .B0(n3564), .B1(n6581), .C0(n7562), 
        .C1(n6617), .Y(N27938) );
  OAI222XL U13245 ( .A0(n7378), .A1(n8014), .B0(n3496), .B1(n8011), .C0(n7562), 
        .C1(n8009), .Y(N28002) );
  OAI222XL U13246 ( .A0(n7378), .A1(n8026), .B0(n3427), .B1(n8024), .C0(n7562), 
        .C1(n8020), .Y(N28066) );
  OAI222XL U13247 ( .A0(n7378), .A1(n8039), .B0(n3359), .B1(n6575), .C0(n7562), 
        .C1(n8033), .Y(N28130) );
  OAI222XL U13248 ( .A0(n7378), .A1(n8079), .B0(n3146), .B1(n8076), .C0(n7562), 
        .C1(n8071), .Y(N28322) );
  OAI222XL U13249 ( .A0(n7378), .A1(n8090), .B0(n3075), .B1(n6578), .C0(n7562), 
        .C1(n8086), .Y(N28386) );
  OAI222XL U13250 ( .A0(n7378), .A1(n8154), .B0(n2592), .B1(n8153), .C0(n7562), 
        .C1(n8150), .Y(N28706) );
  OAI222XL U13251 ( .A0(n7378), .A1(n8169), .B0(n8164), .B1(n2518), .C0(n8162), 
        .C1(n7562), .Y(N28770) );
  AOI221XL U13252 ( .A0(n8764), .A1(n8160), .B0(n8765), .B1(n8146), .C0(n4866), 
        .Y(n4834) );
  CLKINVX1 U13253 ( .A(n2521), .Y(n8764) );
  CLKINVX1 U13254 ( .A(n2593), .Y(n8765) );
  OAI222XL U13255 ( .A0(n8082), .A1(n3076), .B0(n8016), .B1(n3428), .C0(n8069), 
        .C1(n3147), .Y(n4866) );
  AOI221XL U13256 ( .A0(n8759), .A1(n6610), .B0(n8760), .B1(n8144), .C0(n4815), 
        .Y(n4803) );
  CLKINVX1 U13257 ( .A(n2518), .Y(n8759) );
  CLKINVX1 U13258 ( .A(n2592), .Y(n8760) );
  OAI222XL U13259 ( .A0(n8080), .A1(n3075), .B0(n8016), .B1(n3427), .C0(n8068), 
        .C1(n3146), .Y(n4815) );
  OAI221XL U13260 ( .A0(n7376), .A1(n7989), .B0(n7563), .B1(n7986), .C0(n3635), 
        .Y(N27873) );
  OAI221XL U13261 ( .A0(n7376), .A1(n8053), .B0(n7563), .B1(n8050), .C0(n3289), 
        .Y(N28193) );
  OAI221XL U13262 ( .A0(n7376), .A1(n8104), .B0(n7563), .B1(n8101), .C0(n3006), 
        .Y(N28449) );
  OAI221XL U13263 ( .A0(n7376), .A1(n8117), .B0(n7563), .B1(n8114), .C0(n2933), 
        .Y(N28513) );
  OAI221XL U13264 ( .A0(n7376), .A1(n8129), .B0(n7563), .B1(n8127), .C0(n2799), 
        .Y(N28577) );
  OAI221XL U13265 ( .A0(n7376), .A1(n7975), .B0(n7563), .B1(n7973), .C0(n4819), 
        .Y(N27809) );
  OAI221XL U13266 ( .A0(n7378), .A1(n7989), .B0(n7562), .B1(n7986), .C0(n3634), 
        .Y(N27874) );
  OAI221XL U13267 ( .A0(n7378), .A1(n8053), .B0(n7562), .B1(n8050), .C0(n3288), 
        .Y(N28194) );
  OAI221XL U13268 ( .A0(n7378), .A1(n8104), .B0(n7562), .B1(n8101), .C0(n3005), 
        .Y(N28450) );
  OAI221XL U13269 ( .A0(n7378), .A1(n8117), .B0(n7562), .B1(n8114), .C0(n2931), 
        .Y(N28514) );
  OAI221XL U13270 ( .A0(n7378), .A1(n8129), .B0(n7562), .B1(n8127), .C0(n2798), 
        .Y(N28578) );
  OAI221XL U13271 ( .A0(n7378), .A1(n7975), .B0(n7562), .B1(n7973), .C0(n4801), 
        .Y(N27810) );
  CLKINVX1 U13272 ( .A(n3360), .Y(n8767) );
  CLKINVX1 U13273 ( .A(n3359), .Y(n8762) );
  CLKINVX1 U13274 ( .A(n3565), .Y(n8766) );
  CLKINVX1 U13275 ( .A(n3564), .Y(n8761) );
  CLKBUFX3 U13276 ( .A(n8414), .Y(n6990) );
  CLKBUFX3 U13277 ( .A(n8413), .Y(n7002) );
  CLKBUFX3 U13278 ( .A(n8411), .Y(n7007) );
  CLKBUFX3 U13279 ( .A(n6784), .Y(N25537) );
  NAND4X1 U13280 ( .A(n4824), .B(n4825), .C(n4826), .D(n4827), .Y(n3649) );
  NOR4X1 U13281 ( .A(N34888), .B(N34887), .C(N34886), .D(N34885), .Y(n4824) );
  NOR4X1 U13282 ( .A(N34892), .B(N34891), .C(N34890), .D(N34889), .Y(n4825) );
  NOR4BXL U13283 ( .AN(n4831), .B(n4832), .C(n4833), .D(n8883), .Y(n4826) );
  CLKINVX1 U13284 ( .A(N34908), .Y(n8861) );
  NOR4X1 U13285 ( .A(N34908), .B(N34907), .C(N34906), .D(N34905), .Y(n3641) );
  AND4X1 U13286 ( .A(n3640), .B(n3641), .C(n3642), .D(n3643), .Y(n2526) );
  NOR2X1 U13287 ( .A(n3644), .B(n3645), .Y(n3643) );
  NOR4X1 U13288 ( .A(n3648), .B(N34894), .C(N34896), .D(N34895), .Y(n3642) );
  NOR4X1 U13289 ( .A(N34904), .B(N34903), .C(N34902), .D(N34901), .Y(n3640) );
  CLKINVX1 U13290 ( .A(N34903), .Y(n8866) );
  CLKINVX1 U13291 ( .A(N34904), .Y(n8865) );
  CLKINVX1 U13292 ( .A(N34907), .Y(n8862) );
  CLKINVX1 U13293 ( .A(N34906), .Y(n8863) );
  CLKINVX1 U13294 ( .A(N34905), .Y(n8864) );
  CLKINVX1 U13295 ( .A(N34896), .Y(n8873) );
  CLKINVX1 U13296 ( .A(N34902), .Y(n8867) );
  CLKINVX1 U13297 ( .A(N34901), .Y(n8868) );
  CLKINVX1 U13298 ( .A(N34900), .Y(n8869) );
  CLKINVX1 U13299 ( .A(N34899), .Y(n8870) );
  CLKINVX1 U13300 ( .A(N34898), .Y(n8871) );
  CLKINVX1 U13301 ( .A(N34897), .Y(n8872) );
  NOR2BX1 U13302 ( .AN(n4867), .B(n8253), .Y(n4858) );
  NOR2BX1 U13303 ( .AN(n4867), .B(n8184), .Y(n4861) );
  NAND2X1 U13304 ( .A(n4858), .B(n2325), .Y(n3682) );
  NAND4X1 U13305 ( .A(n8878), .B(n8877), .C(n8879), .D(n3647), .Y(n3644) );
  NOR4X1 U13306 ( .A(N34893), .B(N34892), .C(N34891), .D(N34890), .Y(n3647) );
  CLKINVX1 U13307 ( .A(N34895), .Y(n8874) );
  CLKINVX1 U13308 ( .A(N34889), .Y(n8877) );
  CLKINVX1 U13309 ( .A(N34894), .Y(n8875) );
  CLKINVX1 U13310 ( .A(N34893), .Y(n8876) );
  NOR2BX1 U13311 ( .AN(N35114), .B(n8397), .Y(outCount_next[30]) );
  NOR2BX1 U13312 ( .AN(N35113), .B(n8398), .Y(outCount_next[29]) );
  NOR2BX1 U13313 ( .AN(N35112), .B(n159), .Y(outCount_next[28]) );
  NOR2BX1 U13314 ( .AN(N35111), .B(n8397), .Y(outCount_next[27]) );
  AND2X2 U13315 ( .A(N1803), .B(n8405), .Y(N1836) );
  AND2X2 U13316 ( .A(N1802), .B(n8405), .Y(N1835) );
  AND2X2 U13317 ( .A(N1801), .B(n8405), .Y(N1834) );
  AND2X2 U13318 ( .A(N1800), .B(n8405), .Y(N1833) );
  AND2X2 U13319 ( .A(N1799), .B(n8405), .Y(N1832) );
  NAND2X1 U13320 ( .A(n4861), .B(n2325), .Y(n3693) );
  NAND4X1 U13321 ( .A(n241), .B(n8882), .C(n8883), .D(n3646), .Y(n3645) );
  NOR4X1 U13322 ( .A(N34886), .B(N34885), .C(N34884), .D(N34883), .Y(n3646) );
  NAND4X1 U13323 ( .A(n241), .B(n8882), .C(n8881), .D(n8880), .Y(n4832) );
  CLKINVX1 U13324 ( .A(N34882), .Y(n8882) );
  CLKINVX1 U13325 ( .A(N34887), .Y(n8879) );
  CLKINVX1 U13326 ( .A(N34884), .Y(n8880) );
  CLKINVX1 U13327 ( .A(N34888), .Y(n8878) );
  CLKINVX1 U13328 ( .A(N34883), .Y(n8881) );
  NOR2BX1 U13329 ( .AN(N35110), .B(n8397), .Y(outCount_next[26]) );
  NOR2BX1 U13330 ( .AN(N35109), .B(n8397), .Y(outCount_next[25]) );
  NOR2BX1 U13331 ( .AN(N35108), .B(n8397), .Y(outCount_next[24]) );
  NOR2BX1 U13332 ( .AN(N35107), .B(n8397), .Y(outCount_next[23]) );
  NOR2BX1 U13333 ( .AN(N35106), .B(n8397), .Y(outCount_next[22]) );
  NOR2BX1 U13334 ( .AN(N35105), .B(n8397), .Y(outCount_next[21]) );
  NOR2BX1 U13335 ( .AN(N35104), .B(n8397), .Y(outCount_next[20]) );
  AND2X2 U13336 ( .A(N1798), .B(n8405), .Y(N1831) );
  AND2X2 U13337 ( .A(N1797), .B(n8405), .Y(N1830) );
  AND2X2 U13338 ( .A(N1796), .B(n8405), .Y(N1829) );
  AND2X2 U13339 ( .A(N1795), .B(n8405), .Y(N1828) );
  AND2X2 U13340 ( .A(N1794), .B(n8405), .Y(N1827) );
  AND2X2 U13341 ( .A(N1793), .B(n8405), .Y(N1826) );
  AND2X2 U13342 ( .A(N1792), .B(n8405), .Y(N1825) );
  NOR2BX1 U13343 ( .AN(n4867), .B(n8225), .Y(n4849) );
  NOR2BX1 U13344 ( .AN(n4867), .B(n8279), .Y(n4854) );
  NOR2BX1 U13345 ( .AN(n3638), .B(n6988), .Y(n3220) );
  NOR2BX1 U13346 ( .AN(n3078), .B(n6988), .Y(n2523) );
  NOR2BX1 U13347 ( .AN(N35087), .B(n8397), .Y(outCount_next[3]) );
  NOR2BX1 U13348 ( .AN(N35086), .B(n8398), .Y(outCount_next[2]) );
  NAND2X1 U13349 ( .A(n4854), .B(n2325), .Y(n3008) );
  NAND2X1 U13350 ( .A(N34983), .B(n8853), .Y(n135) );
  NAND2X1 U13351 ( .A(n4861), .B(n773), .Y(n2801) );
  NAND2X1 U13352 ( .A(n4849), .B(n2325), .Y(n3291) );
  NAND2X1 U13353 ( .A(n7699), .B(N2348), .Y(n215) );
  NAND2X1 U13354 ( .A(n7687), .B(N2348), .Y(n218) );
  NAND2X1 U13355 ( .A(n7689), .B(N2348), .Y(n222) );
  NAND2X1 U13356 ( .A(n7691), .B(N2348), .Y(n226) );
  NAND2X1 U13357 ( .A(n7693), .B(N2348), .Y(n230) );
  NAND2X1 U13358 ( .A(n7695), .B(N2348), .Y(n234) );
  NAND2X1 U13359 ( .A(n7671), .B(N2348), .Y(n183) );
  NAND2X1 U13360 ( .A(n7673), .B(N2348), .Y(n187) );
  NAND2X1 U13361 ( .A(n7675), .B(N2348), .Y(n191) );
  NAND2X1 U13362 ( .A(n7677), .B(N2348), .Y(n195) );
  NAND2X1 U13363 ( .A(n7679), .B(N2348), .Y(n199) );
  NAND2X1 U13364 ( .A(n7681), .B(N2348), .Y(n203) );
  NAND2X1 U13365 ( .A(n7683), .B(N2348), .Y(n207) );
  NAND2X1 U13366 ( .A(n7685), .B(N2348), .Y(n211) );
  NAND2X1 U13367 ( .A(n7697), .B(N2348), .Y(n238) );
  NAND2X1 U13368 ( .A(N2348), .B(n7669), .Y(n164) );
  CLKINVX1 U13369 ( .A(N34881), .Y(n8883) );
  AND2X2 U13370 ( .A(state_next[0]), .B(state_next[1]), .Y(N35192) );
  CLKBUFX3 U13371 ( .A(n159), .Y(n8397) );
  NOR2BX1 U13372 ( .AN(N34890), .B(n8401), .Y(xCount_next[13]) );
  NOR2BX1 U13373 ( .AN(N34891), .B(n8401), .Y(xCount_next[14]) );
  NOR2BX1 U13374 ( .AN(N34892), .B(n8401), .Y(xCount_next[15]) );
  NOR2BX1 U13375 ( .AN(N35103), .B(n8397), .Y(outCount_next[19]) );
  NOR2BX1 U13376 ( .AN(N35102), .B(n8397), .Y(outCount_next[18]) );
  NOR2BX1 U13377 ( .AN(N35101), .B(n8397), .Y(outCount_next[17]) );
  NOR2BX1 U13378 ( .AN(N35100), .B(n8398), .Y(outCount_next[16]) );
  NOR2BX1 U13379 ( .AN(N35099), .B(n8398), .Y(outCount_next[15]) );
  NOR2BX1 U13380 ( .AN(N35098), .B(n8398), .Y(outCount_next[14]) );
  AND2X2 U13381 ( .A(n3292), .B(n2524), .Y(n181) );
  AND2X2 U13382 ( .A(n2594), .B(n3077), .Y(n189) );
  AND2X2 U13383 ( .A(n2523), .B(n3077), .Y(n193) );
  AND2X2 U13384 ( .A(n2594), .B(n2524), .Y(n213) );
  AND2X2 U13385 ( .A(n3077), .B(n3292), .Y(n4823) );
  AND2X2 U13386 ( .A(n3077), .B(n3220), .Y(n220) );
  AND2X2 U13387 ( .A(n2937), .B(n3292), .Y(n224) );
  AND2X2 U13388 ( .A(n2937), .B(n3220), .Y(n228) );
  AND2X2 U13389 ( .A(n2730), .B(n3292), .Y(n232) );
  AND2X2 U13390 ( .A(n2730), .B(n3220), .Y(n236) );
  AND2X2 U13391 ( .A(n2937), .B(n2594), .Y(n197) );
  AND2X2 U13392 ( .A(n2937), .B(n2523), .Y(n201) );
  AND2X2 U13393 ( .A(n2730), .B(n2594), .Y(n205) );
  AND2X2 U13394 ( .A(n2730), .B(n2523), .Y(n209) );
  CLKBUFX3 U13395 ( .A(n159), .Y(n8398) );
  CLKBUFX3 U13396 ( .A(outCount_next[1]), .Y(n8406) );
  NOR2BX1 U13397 ( .AN(N35085), .B(n8397), .Y(outCount_next[1]) );
  AND2X2 U13398 ( .A(N1791), .B(n8405), .Y(N1824) );
  AND2X2 U13399 ( .A(N1790), .B(n8405), .Y(N1823) );
  AND2X2 U13400 ( .A(N1789), .B(n8405), .Y(N1822) );
  AND2X2 U13401 ( .A(N1788), .B(n8405), .Y(N1821) );
  AND2X2 U13402 ( .A(N1787), .B(n8405), .Y(N1820) );
  AND2X2 U13403 ( .A(N1786), .B(N35189), .Y(N1819) );
  CLKBUFX3 U13404 ( .A(outCount_next[0]), .Y(n7374) );
  CLKINVX1 U13405 ( .A(n161), .Y(n8853) );
  NOR2BX1 U13406 ( .AN(N34885), .B(n8401), .Y(xCount_next[8]) );
  NOR2BX1 U13407 ( .AN(N34886), .B(n8401), .Y(xCount_next[9]) );
  NOR2BX1 U13408 ( .AN(N35093), .B(n159), .Y(outCount_next[9]) );
  NOR2BX1 U13409 ( .AN(N35092), .B(n159), .Y(outCount_next[8]) );
  NOR2BX1 U13410 ( .AN(N35091), .B(n159), .Y(outCount_next[7]) );
  NOR2BX1 U13411 ( .AN(N35090), .B(n8397), .Y(outCount_next[6]) );
  NOR2BX1 U13412 ( .AN(N35089), .B(n8398), .Y(outCount_next[5]) );
  NOR2BX1 U13413 ( .AN(N35088), .B(n8397), .Y(outCount_next[4]) );
  NOR2BX1 U13414 ( .AN(N35097), .B(n8398), .Y(outCount_next[13]) );
  NOR2BX1 U13415 ( .AN(N35096), .B(n8398), .Y(outCount_next[12]) );
  NOR2BX1 U13416 ( .AN(N35095), .B(n8398), .Y(outCount_next[11]) );
  NOR2BX1 U13417 ( .AN(N35094), .B(n8398), .Y(outCount_next[10]) );
  OAI2BB1X1 U13418 ( .A0N(N1777), .A1N(n8405), .B0(n4883), .Y(N1810) );
  AND2X2 U13419 ( .A(N1785), .B(N35189), .Y(N1818) );
  AND2X2 U13420 ( .A(N1784), .B(N35189), .Y(N1817) );
  AND2X2 U13421 ( .A(N1783), .B(N35189), .Y(N1816) );
  AND2X2 U13422 ( .A(N1782), .B(N35189), .Y(N1815) );
  AND2X2 U13423 ( .A(N1781), .B(N35189), .Y(N1814) );
  AND2X2 U13424 ( .A(N1780), .B(N35189), .Y(N1813) );
  AND2X2 U13425 ( .A(N1779), .B(N35189), .Y(N1812) );
  AND2X2 U13426 ( .A(N1774), .B(n8404), .Y(N1807) );
  AND2X2 U13427 ( .A(N1773), .B(n8404), .Y(N1806) );
  AND2X2 U13428 ( .A(N1778), .B(N35189), .Y(N1811) );
  AND2X2 U13429 ( .A(N1776), .B(N35189), .Y(N1809) );
  AND2X2 U13430 ( .A(N1775), .B(N35189), .Y(N1808) );
  OAI221XL U13431 ( .A0(n8315), .A1(n271), .B0(n7737), .B1(n267), .C0(n783), 
        .Y(N34025) );
  OAI221XL U13432 ( .A0(n8312), .A1(n1296), .B0(n7714), .B1(n1298), .C0(n1552), 
        .Y(N33833) );
  CLKBUFX3 U13433 ( .A(n8830), .Y(n7569) );
  CLKBUFX3 U13434 ( .A(n8830), .Y(n7568) );
  CLKBUFX3 U13435 ( .A(n8830), .Y(n7567) );
  OAI221X1 U13436 ( .A0(\xArray[7][1] ), .A1(n8295), .B0(\xArray[11][1] ), 
        .B1(n8241), .C0(n1289), .Y(n765) );
  AOI2BB2X1 U13437 ( .B0(n9384), .B1(n8210), .A0N(\xArray[15][1] ), .A1N(n8254), .Y(n1289) );
  OA22X1 U13438 ( .A0(\xArray[0][3] ), .A1(n8189), .B0(\xArray[12][3] ), .B1(
        n8261), .Y(n2296) );
  OA22X1 U13439 ( .A0(\xArray[0][4] ), .A1(n8189), .B0(\xArray[12][4] ), .B1(
        n8262), .Y(n2287) );
  OAI221X1 U13440 ( .A0(\xArray[8][1] ), .A1(n8295), .B0(\xArray[12][1] ), 
        .B1(n8241), .C0(n1288), .Y(n767) );
  OA22X1 U13441 ( .A0(\xArray[4][1] ), .A1(n8198), .B0(\xArray[0][1] ), .B1(
        n8270), .Y(n1288) );
  OAI221X1 U13442 ( .A0(\xArray[6][1] ), .A1(n8292), .B0(\xArray[10][1] ), 
        .B1(n8238), .C0(n1547), .Y(n971) );
  OAI221X1 U13443 ( .A0(\xArray[6][2] ), .A1(n8292), .B0(\xArray[10][2] ), 
        .B1(n8238), .C0(n1543), .Y(n968) );
  OAI221X1 U13444 ( .A0(\xArray[6][3] ), .A1(n8292), .B0(\xArray[10][3] ), 
        .B1(n8238), .C0(n1539), .Y(n965) );
  OA22X1 U13445 ( .A0(\xArray[14][3] ), .A1(n8273), .B0(\xArray[2][3] ), .B1(
        n8187), .Y(n1539) );
  OA22X1 U13446 ( .A0(\xArray[1][4] ), .A1(n8187), .B0(\xArray[13][4] ), .B1(
        n8260), .Y(n1731) );
  OAI221X1 U13447 ( .A0(\xArray[5][1] ), .A1(n8280), .B0(\xArray[9][1] ), .B1(
        n8226), .C0(n1740), .Y(n1287) );
  OAI221XL U13448 ( .A0(\xArray[9][1] ), .A1(n8290), .B0(\xArray[13][1] ), 
        .B1(n8236), .C0(n972), .Y(n766) );
  OA22X1 U13449 ( .A0(\xArray[5][1] ), .A1(n8196), .B0(\xArray[1][1] ), .B1(
        n8268), .Y(n972) );
  OAI221XL U13450 ( .A0(n7487), .A1(n8065), .B0(n7507), .B1(n8063), .C0(n3161), 
        .Y(N28313) );
  OAI221XL U13451 ( .A0(n7487), .A1(n8143), .B0(n7507), .B1(n8140), .C0(n2614), 
        .Y(N28697) );
  OAI221XL U13452 ( .A0(n7489), .A1(n8066), .B0(n7506), .B1(n8063), .C0(n3160), 
        .Y(N28314) );
  OAI221XL U13453 ( .A0(n7489), .A1(n8143), .B0(n7506), .B1(n8140), .C0(n2612), 
        .Y(N28698) );
  OAI221XL U13454 ( .A0(n7491), .A1(n8065), .B0(n7505), .B1(n8062), .C0(n3159), 
        .Y(N28315) );
  OAI221XL U13455 ( .A0(n7491), .A1(n6608), .B0(n7505), .B1(n8139), .C0(n2610), 
        .Y(N28699) );
  OAI221XL U13456 ( .A0(n7493), .A1(n8065), .B0(n7504), .B1(n8061), .C0(n3158), 
        .Y(N28316) );
  OAI221XL U13457 ( .A0(n7493), .A1(n8142), .B0(n7504), .B1(n8138), .C0(n2608), 
        .Y(N28700) );
  OAI221XL U13458 ( .A0(n7495), .A1(n8065), .B0(n7503), .B1(n6593), .C0(n3157), 
        .Y(N28317) );
  OAI221XL U13459 ( .A0(n7495), .A1(n8142), .B0(n7503), .B1(n6594), .C0(n2606), 
        .Y(N28701) );
  OAI221XL U13460 ( .A0(n7497), .A1(n6607), .B0(n7566), .B1(n6593), .C0(n3156), 
        .Y(N28318) );
  OAI221XL U13461 ( .A0(n7497), .A1(n8142), .B0(n7566), .B1(n6594), .C0(n2604), 
        .Y(N28702) );
  OAI221XL U13462 ( .A0(n7499), .A1(n8066), .B0(n7566), .B1(n6593), .C0(n3155), 
        .Y(N28319) );
  OAI221XL U13463 ( .A0(n7499), .A1(n8143), .B0(n7566), .B1(n6594), .C0(n2602), 
        .Y(N28703) );
  OAI221XL U13464 ( .A0(n7501), .A1(n6607), .B0(n7566), .B1(n6593), .C0(n3152), 
        .Y(N28320) );
  OAI221XL U13465 ( .A0(n7501), .A1(n6608), .B0(n7565), .B1(n6594), .C0(n2598), 
        .Y(N28704) );
  OAI22X1 U13466 ( .A0(\xArray[0][57] ), .A1(n7770), .B0(n7777), .B1(n7488), 
        .Y(n2350) );
  OAI22X1 U13467 ( .A0(\xArray[0][58] ), .A1(n7770), .B0(n7776), .B1(n7490), 
        .Y(n2347) );
  OAI22X1 U13468 ( .A0(\xArray[0][59] ), .A1(n7771), .B0(n7776), .B1(n7492), 
        .Y(n2344) );
  OAI22X1 U13469 ( .A0(\xArray[0][60] ), .A1(n7773), .B0(n7775), .B1(n7494), 
        .Y(n2341) );
  OAI22X1 U13470 ( .A0(\xArray[0][61] ), .A1(n7773), .B0(n7775), .B1(n7496), 
        .Y(n2338) );
  OAI22X1 U13471 ( .A0(\xArray[0][62] ), .A1(n7771), .B0(n7774), .B1(n7498), 
        .Y(n2335) );
  OAI22X1 U13472 ( .A0(\xArray[0][63] ), .A1(n7768), .B0(n7774), .B1(n7500), 
        .Y(n2331) );
  OAI22X1 U13473 ( .A0(\xArray[1][57] ), .A1(n7785), .B0(n7801), .B1(n7488), 
        .Y(n2536) );
  OAI22X1 U13474 ( .A0(\xArray[1][58] ), .A1(n7785), .B0(n7799), .B1(n7490), 
        .Y(n2535) );
  OAI22X1 U13475 ( .A0(\xArray[1][59] ), .A1(n7785), .B0(n7798), .B1(n7492), 
        .Y(n2534) );
  OAI22X1 U13476 ( .A0(\xArray[1][60] ), .A1(n7785), .B0(n7797), .B1(n7494), 
        .Y(n2533) );
  OAI22X1 U13477 ( .A0(\xArray[10][60] ), .A1(n7890), .B0(n7907), .B1(n7494), 
        .Y(n3300) );
  OAI22X1 U13478 ( .A0(\xArray[13][60] ), .A1(n7871), .B0(n7879), .B1(n7494), 
        .Y(n3505) );
  OAI22X1 U13479 ( .A0(\xArray[1][61] ), .A1(n7785), .B0(n7796), .B1(n7496), 
        .Y(n2532) );
  OAI22X1 U13480 ( .A0(\xArray[1][62] ), .A1(n7785), .B0(n7795), .B1(n7498), 
        .Y(n2531) );
  OAI22X1 U13481 ( .A0(\xArray[1][63] ), .A1(n7785), .B0(n7794), .B1(n7500), 
        .Y(n2528) );
  OAI22X1 U13482 ( .A0(\xArray[13][63] ), .A1(n7868), .B0(n7876), .B1(n7500), 
        .Y(n3500) );
  OAI22X1 U13483 ( .A0(\xArray[10][63] ), .A1(n7890), .B0(n7500), .B1(n7902), 
        .Y(n3295) );
  OAI22X1 U13484 ( .A0(\xArray[7][56] ), .A1(n7850), .B0(n7863), .B1(n7486), 
        .Y(n3091) );
  OAI22X1 U13485 ( .A0(\xArray[7][57] ), .A1(n7850), .B0(n7863), .B1(n7488), 
        .Y(n3090) );
  OAI22X1 U13486 ( .A0(\xArray[7][58] ), .A1(n7850), .B0(n7864), .B1(n7490), 
        .Y(n3089) );
  OAI22X1 U13487 ( .A0(\xArray[7][59] ), .A1(n7850), .B0(n7864), .B1(n7492), 
        .Y(n3088) );
  OAI22X1 U13488 ( .A0(\xArray[7][60] ), .A1(n7848), .B0(n7864), .B1(n7494), 
        .Y(n3087) );
  OAI22X1 U13489 ( .A0(\xArray[12][60] ), .A1(n7909), .B0(n7925), .B1(n7494), 
        .Y(n3437) );
  OAI22X1 U13490 ( .A0(\xArray[7][61] ), .A1(n7848), .B0(n7864), .B1(n7496), 
        .Y(n3086) );
  OAI22X1 U13491 ( .A0(\xArray[7][62] ), .A1(n7848), .B0(n7865), .B1(n7498), 
        .Y(n3085) );
  OAI22X1 U13492 ( .A0(\xArray[6][56] ), .A1(n7809), .B0(n7821), .B1(n7486), 
        .Y(n3020) );
  OAI22X1 U13493 ( .A0(\xArray[6][57] ), .A1(n7809), .B0(n7821), .B1(n7488), 
        .Y(n3019) );
  OAI22X1 U13494 ( .A0(\xArray[6][58] ), .A1(n7809), .B0(n7822), .B1(n7490), 
        .Y(n3018) );
  OAI22X1 U13495 ( .A0(\xArray[6][59] ), .A1(n7809), .B0(n7822), .B1(n7492), 
        .Y(n3017) );
  OAI22X1 U13496 ( .A0(\xArray[6][60] ), .A1(n7809), .B0(n7822), .B1(n7494), 
        .Y(n3016) );
  OAI22X1 U13497 ( .A0(\xArray[6][61] ), .A1(n7810), .B0(n7822), .B1(n7496), 
        .Y(n3015) );
  OAI22X1 U13498 ( .A0(\xArray[6][62] ), .A1(n7808), .B0(n7823), .B1(n7498), 
        .Y(n3014) );
  OAI22X1 U13499 ( .A0(\xArray[11][56] ), .A1(n7828), .B0(n7843), .B1(n7486), 
        .Y(n3372) );
  OAI22X1 U13500 ( .A0(\xArray[11][57] ), .A1(n7828), .B0(n7843), .B1(n7488), 
        .Y(n3371) );
  OAI22X1 U13501 ( .A0(\xArray[11][58] ), .A1(n7828), .B0(n7841), .B1(n7490), 
        .Y(n3370) );
  OAI22X1 U13502 ( .A0(\xArray[11][59] ), .A1(n7828), .B0(n7842), .B1(n7492), 
        .Y(n3369) );
  OAI22X1 U13503 ( .A0(\xArray[11][60] ), .A1(n7829), .B0(n7844), .B1(n7494), 
        .Y(n3368) );
  OAI22X1 U13504 ( .A0(\xArray[11][61] ), .A1(n7829), .B0(n7841), .B1(n7496), 
        .Y(n3367) );
  OAI22X1 U13505 ( .A0(\xArray[11][62] ), .A1(n7829), .B0(n7844), .B1(n7498), 
        .Y(n3366) );
  OAI22X1 U13506 ( .A0(\xArray[7][63] ), .A1(n7848), .B0(n7500), .B1(n7865), 
        .Y(n3082) );
  OAI22X1 U13507 ( .A0(\xArray[12][63] ), .A1(n7909), .B0(n7500), .B1(n7925), 
        .Y(n3432) );
  OAI22X1 U13508 ( .A0(\xArray[6][63] ), .A1(n7810), .B0(n7500), .B1(n7823), 
        .Y(n3011) );
  OAI22X1 U13509 ( .A0(\xArray[11][63] ), .A1(n7829), .B0(n7500), .B1(n7844), 
        .Y(n3363) );
  AND4X1 U13510 ( .A(n3813), .B(n3814), .C(n3815), .D(n3816), .Y(n2352) );
  AOI221XL U13511 ( .A0(n7963), .A1(\xArray[9][56] ), .B0(\xArray[8][56] ), 
        .B1(n7959), .C0(n3817), .Y(n3816) );
  AOI221XL U13512 ( .A0(n7947), .A1(n7486), .B0(n3667), .B1(\xArray[2][56] ), 
        .C0(n3819), .Y(n3815) );
  AND4X1 U13513 ( .A(n3795), .B(n3796), .C(n3797), .D(n3798), .Y(n2349) );
  AOI221XL U13514 ( .A0(n7963), .A1(\xArray[9][57] ), .B0(\xArray[8][57] ), 
        .B1(n7959), .C0(n3799), .Y(n3798) );
  AOI221XL U13515 ( .A0(n7947), .A1(n7488), .B0(n7946), .B1(\xArray[2][57] ), 
        .C0(n3801), .Y(n3797) );
  AND4X1 U13516 ( .A(n3777), .B(n3778), .C(n3779), .D(n3780), .Y(n2346) );
  AOI221XL U13517 ( .A0(n7963), .A1(\xArray[9][58] ), .B0(\xArray[8][58] ), 
        .B1(n7959), .C0(n3781), .Y(n3780) );
  AOI221XL U13518 ( .A0(n7947), .A1(n7490), .B0(n7945), .B1(\xArray[2][58] ), 
        .C0(n3783), .Y(n3779) );
  AND4X1 U13519 ( .A(n3759), .B(n3760), .C(n3761), .D(n3762), .Y(n2343) );
  AOI221XL U13520 ( .A0(n7963), .A1(\xArray[9][59] ), .B0(\xArray[8][59] ), 
        .B1(n7959), .C0(n3763), .Y(n3762) );
  AOI221XL U13521 ( .A0(n7947), .A1(n7492), .B0(n3667), .B1(\xArray[2][59] ), 
        .C0(n3765), .Y(n3761) );
  BUFX4 U13522 ( .A(n2340), .Y(n7495) );
  AND4X1 U13523 ( .A(n3741), .B(n3742), .C(n3743), .D(n3744), .Y(n2340) );
  AOI221XL U13524 ( .A0(n7963), .A1(\xArray[9][60] ), .B0(\xArray[8][60] ), 
        .B1(n7959), .C0(n3745), .Y(n3744) );
  AOI221XL U13525 ( .A0(n7947), .A1(n7494), .B0(n7946), .B1(\xArray[2][60] ), 
        .C0(n3747), .Y(n3743) );
  AND4X1 U13526 ( .A(n3723), .B(n3724), .C(n3725), .D(n3726), .Y(n2337) );
  AOI221XL U13527 ( .A0(n7963), .A1(\xArray[9][61] ), .B0(\xArray[8][61] ), 
        .B1(n7959), .C0(n3727), .Y(n3726) );
  AOI221XL U13528 ( .A0(n7947), .A1(n7496), .B0(n7945), .B1(\xArray[2][61] ), 
        .C0(n3729), .Y(n3725) );
  AND4X1 U13529 ( .A(n3705), .B(n3706), .C(n3707), .D(n3708), .Y(n2334) );
  AOI221XL U13530 ( .A0(n7963), .A1(\xArray[9][62] ), .B0(\xArray[8][62] ), 
        .B1(n7959), .C0(n3709), .Y(n3708) );
  AOI221XL U13531 ( .A0(n7947), .A1(n7498), .B0(n7946), .B1(\xArray[2][62] ), 
        .C0(n3711), .Y(n3707) );
  AND4X1 U13532 ( .A(n3655), .B(n3656), .C(n3657), .D(n3658), .Y(n2328) );
  AOI221XL U13533 ( .A0(n7963), .A1(\xArray[9][63] ), .B0(\xArray[8][63] ), 
        .B1(n7959), .C0(n3661), .Y(n3658) );
  AOI221XL U13534 ( .A0(n7947), .A1(n7500), .B0(n7945), .B1(\xArray[2][63] ), 
        .C0(n3668), .Y(n3657) );
  OAI221X1 U13535 ( .A0(\xArray[7][2] ), .A1(n8295), .B0(\xArray[11][2] ), 
        .B1(n8241), .C0(n1284), .Y(n757) );
  AOI2BB2X1 U13536 ( .B0(n9376), .B1(n8210), .A0N(\xArray[15][2] ), .A1N(n8254), .Y(n1284) );
  OAI221X1 U13537 ( .A0(\xArray[7][3] ), .A1(n8295), .B0(\xArray[11][3] ), 
        .B1(n8241), .C0(n1279), .Y(n749) );
  OA22X1 U13538 ( .A0(\xArray[0][2] ), .A1(n8189), .B0(\xArray[12][2] ), .B1(
        n8261), .Y(n2305) );
  OA22X1 U13539 ( .A0(\xArray[0][5] ), .A1(n8189), .B0(\xArray[12][5] ), .B1(
        n8262), .Y(n2278) );
  OAI221X1 U13540 ( .A0(\xArray[4][6] ), .A1(n8284), .B0(\xArray[8][6] ), .B1(
        n8230), .C0(n2269), .Y(n1524) );
  OA22X1 U13541 ( .A0(\xArray[4][2] ), .A1(n8198), .B0(\xArray[0][2] ), .B1(
        n8270), .Y(n1283) );
  OAI221X1 U13542 ( .A0(\xArray[8][3] ), .A1(n8295), .B0(\xArray[12][3] ), 
        .B1(n8241), .C0(n1278), .Y(n751) );
  OAI221X1 U13543 ( .A0(\xArray[8][4] ), .A1(n8295), .B0(\xArray[12][4] ), 
        .B1(n8241), .C0(n1273), .Y(n743) );
  OAI221X1 U13544 ( .A0(\xArray[8][5] ), .A1(n8295), .B0(\xArray[12][5] ), 
        .B1(n8241), .C0(n1268), .Y(n735) );
  OA22X1 U13545 ( .A0(\xArray[15][3] ), .A1(n8189), .B0(\xArray[11][3] ), .B1(
        n8262), .Y(n2295) );
  OAI221X1 U13546 ( .A0(\xArray[3][4] ), .A1(n8283), .B0(\xArray[7][4] ), .B1(
        n8229), .C0(n2286), .Y(n1534) );
  OA22X1 U13547 ( .A0(\xArray[15][4] ), .A1(n8189), .B0(\xArray[11][4] ), .B1(
        n8262), .Y(n2286) );
  OAI221X1 U13548 ( .A0(\xArray[3][5] ), .A1(n8284), .B0(\xArray[7][5] ), .B1(
        n8230), .C0(n2277), .Y(n1530) );
  OA22X1 U13549 ( .A0(\xArray[15][5] ), .A1(n8189), .B0(\xArray[11][5] ), .B1(
        n8263), .Y(n2277) );
  OA22X1 U13550 ( .A0(\xArray[14][0] ), .A1(n8272), .B0(\xArray[2][0] ), .B1(
        n8187), .Y(n1551) );
  OA22X1 U13551 ( .A0(\xArray[1][3] ), .A1(n8187), .B0(\xArray[13][3] ), .B1(
        n8260), .Y(n1734) );
  OAI221X1 U13552 ( .A0(\xArray[5][5] ), .A1(n8281), .B0(\xArray[9][5] ), .B1(
        n8227), .C0(n1728), .Y(n1267) );
  OA22X1 U13553 ( .A0(\xArray[1][5] ), .A1(n8187), .B0(\xArray[13][5] ), .B1(
        n8260), .Y(n1728) );
  AOI2BB2X1 U13554 ( .B0(n9392), .B1(n8210), .A0N(\xArray[15][0] ), .A1N(n8254), .Y(n1294) );
  OAI221X1 U13555 ( .A0(\xArray[8][0] ), .A1(n8295), .B0(\xArray[12][0] ), 
        .B1(n8241), .C0(n1293), .Y(n782) );
  OA22X1 U13556 ( .A0(\xArray[4][0] ), .A1(n8198), .B0(\xArray[0][0] ), .B1(
        n8270), .Y(n1293) );
  OAI221X1 U13557 ( .A0(\xArray[5][0] ), .A1(n8280), .B0(\xArray[9][0] ), .B1(
        n8226), .C0(n1743), .Y(n1292) );
  OA22X1 U13558 ( .A0(\xArray[1][0] ), .A1(n8187), .B0(\xArray[13][0] ), .B1(
        n8260), .Y(n1743) );
  OAI221X1 U13559 ( .A0(\xArray[3][0] ), .A1(n8283), .B0(\xArray[7][0] ), .B1(
        n8229), .C0(n2326), .Y(n1550) );
  OAI221XL U13560 ( .A0(\xArray[9][3] ), .A1(n8290), .B0(\xArray[13][3] ), 
        .B1(n8236), .C0(n966), .Y(n750) );
  OA22X1 U13561 ( .A0(\xArray[5][3] ), .A1(n8196), .B0(\xArray[1][3] ), .B1(
        n8268), .Y(n966) );
  OAI221XL U13562 ( .A0(\xArray[9][4] ), .A1(n8290), .B0(\xArray[13][4] ), 
        .B1(n8236), .C0(n963), .Y(n742) );
  OA22X1 U13563 ( .A0(\xArray[5][0] ), .A1(n8196), .B0(\xArray[1][0] ), .B1(
        n8268), .Y(n975) );
  OAI221XL U13564 ( .A0(\xArray[2][1] ), .A1(n8283), .B0(\xArray[6][1] ), .B1(
        n8229), .C0(n2311), .Y(n1739) );
  AOI221XL U13565 ( .A0(n7947), .A1(n7478), .B0(n7944), .B1(\xArray[2][52] ), 
        .C0(n3891), .Y(n3887) );
  OAI222XL U13566 ( .A0(n8978), .A1(n7941), .B0(n8503), .B1(n7938), .C0(n7936), 
        .C1(n8977), .Y(n3891) );
  OAI221XL U13567 ( .A0(n7479), .A1(n6607), .B0(n7511), .B1(n6593), .C0(n3165), 
        .Y(N28309) );
  OAI221XL U13568 ( .A0(n7479), .A1(n6608), .B0(n7511), .B1(n6594), .C0(n2622), 
        .Y(N28693) );
  OAI221XL U13569 ( .A0(n7481), .A1(n8064), .B0(n7510), .B1(n6593), .C0(n3164), 
        .Y(N28310) );
  OAI221XL U13570 ( .A0(n7481), .A1(n8141), .B0(n7510), .B1(n6594), .C0(n2620), 
        .Y(N28694) );
  OAI221XL U13571 ( .A0(n7483), .A1(n8065), .B0(n7509), .B1(n8061), .C0(n3163), 
        .Y(N28311) );
  OAI221XL U13572 ( .A0(n7483), .A1(n8142), .B0(n7509), .B1(n8138), .C0(n2618), 
        .Y(N28695) );
  OAI221XL U13573 ( .A0(n7485), .A1(n8065), .B0(n7508), .B1(n8061), .C0(n3162), 
        .Y(N28312) );
  OAI221XL U13574 ( .A0(n7485), .A1(n8142), .B0(n7508), .B1(n8138), .C0(n2616), 
        .Y(N28696) );
  OAI22X1 U13575 ( .A0(\xArray[0][55] ), .A1(n7771), .B0(n7778), .B1(n7484), 
        .Y(n2356) );
  OAI22X1 U13576 ( .A0(\xArray[0][56] ), .A1(n7771), .B0(n7777), .B1(n7486), 
        .Y(n2353) );
  OAI22X1 U13577 ( .A0(\xArray[1][55] ), .A1(n7786), .B0(n7802), .B1(n7484), 
        .Y(n2538) );
  OAI22X1 U13578 ( .A0(\xArray[1][56] ), .A1(n7785), .B0(n7799), .B1(n7486), 
        .Y(n2537) );
  OAI22X1 U13579 ( .A0(\xArray[7][53] ), .A1(n7850), .B0(n7861), .B1(n7480), 
        .Y(n3094) );
  OAI22X1 U13580 ( .A0(\xArray[7][54] ), .A1(n7850), .B0(n7863), .B1(n7482), 
        .Y(n3093) );
  OAI22X1 U13581 ( .A0(\xArray[7][55] ), .A1(n7848), .B0(n7863), .B1(n7484), 
        .Y(n3092) );
  OAI22X1 U13582 ( .A0(\xArray[6][53] ), .A1(n7809), .B0(n7822), .B1(n7480), 
        .Y(n3023) );
  OAI22X1 U13583 ( .A0(\xArray[6][54] ), .A1(n7810), .B0(n7821), .B1(n7482), 
        .Y(n3022) );
  OAI22X1 U13584 ( .A0(\xArray[6][55] ), .A1(n7810), .B0(n7821), .B1(n7484), 
        .Y(n3021) );
  OAI22X1 U13585 ( .A0(\xArray[11][55] ), .A1(n7829), .B0(n7843), .B1(n7484), 
        .Y(n3373) );
  AND4X1 U13586 ( .A(n3867), .B(n3868), .C(n3869), .D(n3870), .Y(n2361) );
  AOI221XL U13587 ( .A0(n7963), .A1(\xArray[9][53] ), .B0(\xArray[8][53] ), 
        .B1(n7959), .C0(n3871), .Y(n3870) );
  AOI221XL U13588 ( .A0(n7947), .A1(n7480), .B0(n7946), .B1(\xArray[2][53] ), 
        .C0(n3873), .Y(n3869) );
  AND4X1 U13589 ( .A(n3849), .B(n3850), .C(n3851), .D(n3852), .Y(n2358) );
  AOI221XL U13590 ( .A0(n7963), .A1(\xArray[9][54] ), .B0(\xArray[8][54] ), 
        .B1(n7959), .C0(n3853), .Y(n3852) );
  AOI221XL U13591 ( .A0(n7947), .A1(n7482), .B0(n7945), .B1(\xArray[2][54] ), 
        .C0(n3855), .Y(n3851) );
  AND4X1 U13592 ( .A(n3831), .B(n3832), .C(n3833), .D(n3834), .Y(n2355) );
  AOI221XL U13593 ( .A0(n7963), .A1(\xArray[9][55] ), .B0(\xArray[8][55] ), 
        .B1(n7959), .C0(n3835), .Y(n3834) );
  AOI221XL U13594 ( .A0(n7947), .A1(n7484), .B0(n7944), .B1(\xArray[2][55] ), 
        .C0(n3837), .Y(n3833) );
  OAI221X1 U13595 ( .A0(\xArray[4][7] ), .A1(n8284), .B0(\xArray[8][7] ), .B1(
        n8230), .C0(n2260), .Y(n1520) );
  OAI221X1 U13596 ( .A0(\xArray[8][6] ), .A1(n8295), .B0(\xArray[12][6] ), 
        .B1(n8241), .C0(n1263), .Y(n727) );
  OAI221X1 U13597 ( .A0(\xArray[6][6] ), .A1(n8292), .B0(\xArray[10][6] ), 
        .B1(n8238), .C0(n1527), .Y(n956) );
  OAI221X1 U13598 ( .A0(\xArray[3][6] ), .A1(n8284), .B0(\xArray[7][6] ), .B1(
        n8230), .C0(n2268), .Y(n1526) );
  OAI221X1 U13599 ( .A0(\xArray[6][7] ), .A1(n8292), .B0(\xArray[10][7] ), 
        .B1(n8238), .C0(n1523), .Y(n953) );
  OAI221X1 U13600 ( .A0(\xArray[3][7] ), .A1(n8284), .B0(\xArray[7][7] ), .B1(
        n8230), .C0(n2259), .Y(n1522) );
  OAI221X1 U13601 ( .A0(\xArray[5][7] ), .A1(n8281), .B0(\xArray[9][7] ), .B1(
        n8227), .C0(n1722), .Y(n1257) );
  OAI221X1 U13602 ( .A0(\xArray[4][0] ), .A1(n8286), .B0(\xArray[8][0] ), .B1(
        n8232), .C0(n2327), .Y(n1548) );
  OA22X1 U13603 ( .A0(\xArray[0][0] ), .A1(n8192), .B0(\xArray[12][0] ), .B1(
        n8260), .Y(n2327) );
  OAI221XL U13604 ( .A0(\xArray[9][5] ), .A1(n8290), .B0(\xArray[13][5] ), 
        .B1(n8236), .C0(n960), .Y(n734) );
  OAI221XL U13605 ( .A0(\xArray[9][6] ), .A1(n8290), .B0(\xArray[13][6] ), 
        .B1(n8236), .C0(n957), .Y(n726) );
  OAI221XL U13606 ( .A0(\xArray[2][3] ), .A1(n8283), .B0(\xArray[6][3] ), .B1(
        n8229), .C0(n2293), .Y(n1733) );
  AOI2BB2X1 U13607 ( .B0(n9374), .B1(n8207), .A0N(\xArray[10][3] ), .A1N(n8257), .Y(n2293) );
  OAI221XL U13608 ( .A0(\xArray[2][4] ), .A1(n8283), .B0(\xArray[6][4] ), .B1(
        n8229), .C0(n2284), .Y(n1730) );
  AOI2BB2X1 U13609 ( .B0(n9366), .B1(n8207), .A0N(\xArray[10][4] ), .A1N(n8257), .Y(n2284) );
  AOI2BB2X1 U13610 ( .B0(n9398), .B1(n8210), .A0N(\xArray[10][0] ), .A1N(n8258), .Y(n2323) );
  AOI221XL U13611 ( .A0(n7948), .A1(n7476), .B0(n7945), .B1(\xArray[2][51] ), 
        .C0(n3909), .Y(n3905) );
  OAI222XL U13612 ( .A0(n8986), .A1(n7942), .B0(n8508), .B1(n7939), .C0(n7936), 
        .C1(n8985), .Y(n3909) );
  OAI221XL U13613 ( .A0(n7473), .A1(n8066), .B0(n7514), .B1(n8063), .C0(n3168), 
        .Y(N28306) );
  OAI221XL U13614 ( .A0(n7473), .A1(n8142), .B0(n7514), .B1(n8140), .C0(n2628), 
        .Y(N28690) );
  OAI221XL U13615 ( .A0(n7475), .A1(n8066), .B0(n7513), .B1(n8063), .C0(n3167), 
        .Y(N28307) );
  OAI221XL U13616 ( .A0(n7475), .A1(n8143), .B0(n7513), .B1(n8140), .C0(n2626), 
        .Y(N28691) );
  OAI221XL U13617 ( .A0(n7477), .A1(n8064), .B0(n7512), .B1(n8061), .C0(n3166), 
        .Y(N28308) );
  OAI221XL U13618 ( .A0(n7477), .A1(n8141), .B0(n7512), .B1(n8138), .C0(n2624), 
        .Y(N28692) );
  OAI22X1 U13619 ( .A0(\xArray[7][49] ), .A1(n7849), .B0(n7862), .B1(n7472), 
        .Y(n3098) );
  OAI22X1 U13620 ( .A0(\xArray[7][50] ), .A1(n7849), .B0(n7864), .B1(n7474), 
        .Y(n3097) );
  OAI22X1 U13621 ( .A0(\xArray[6][49] ), .A1(n7808), .B0(n7821), .B1(n7472), 
        .Y(n3027) );
  OAI22X1 U13622 ( .A0(\xArray[6][50] ), .A1(n7808), .B0(n7821), .B1(n7474), 
        .Y(n3026) );
  AND4X1 U13623 ( .A(n3939), .B(n3940), .C(n3941), .D(n3942), .Y(n2373) );
  AOI221XL U13624 ( .A0(n7964), .A1(\xArray[9][49] ), .B0(\xArray[8][49] ), 
        .B1(n7960), .C0(n3943), .Y(n3942) );
  AOI221XL U13625 ( .A0(n7948), .A1(n7472), .B0(n7945), .B1(\xArray[2][49] ), 
        .C0(n3945), .Y(n3941) );
  AND4X1 U13626 ( .A(n3921), .B(n3922), .C(n3923), .D(n3924), .Y(n2370) );
  AOI221XL U13627 ( .A0(n7964), .A1(\xArray[9][50] ), .B0(\xArray[8][50] ), 
        .B1(n7960), .C0(n3925), .Y(n3924) );
  AOI221XL U13628 ( .A0(n7948), .A1(n7474), .B0(n7945), .B1(\xArray[2][50] ), 
        .C0(n3927), .Y(n3923) );
  OAI221X1 U13629 ( .A0(\xArray[7][9] ), .A1(n8296), .B0(\xArray[11][9] ), 
        .B1(n8242), .C0(n1249), .Y(n701) );
  OAI221X1 U13630 ( .A0(\xArray[4][9] ), .A1(n8284), .B0(\xArray[8][9] ), .B1(
        n8230), .C0(n2242), .Y(n1512) );
  OA22X1 U13631 ( .A0(\xArray[0][9] ), .A1(n8190), .B0(\xArray[12][9] ), .B1(
        n8264), .Y(n2242) );
  OAI221X1 U13632 ( .A0(\xArray[8][7] ), .A1(n8295), .B0(\xArray[12][7] ), 
        .B1(n8241), .C0(n1258), .Y(n719) );
  OAI221X1 U13633 ( .A0(\xArray[8][8] ), .A1(n8296), .B0(\xArray[12][8] ), 
        .B1(n8242), .C0(n1253), .Y(n711) );
  OA22X1 U13634 ( .A0(\xArray[4][8] ), .A1(n8198), .B0(\xArray[0][8] ), .B1(
        n8270), .Y(n1253) );
  OAI221X1 U13635 ( .A0(\xArray[6][8] ), .A1(n8292), .B0(\xArray[10][8] ), 
        .B1(n8238), .C0(n1519), .Y(n950) );
  OAI221X1 U13636 ( .A0(\xArray[3][8] ), .A1(n8284), .B0(\xArray[7][8] ), .B1(
        n8230), .C0(n2250), .Y(n1518) );
  OAI221X1 U13637 ( .A0(\xArray[6][9] ), .A1(n8292), .B0(\xArray[10][9] ), 
        .B1(n8238), .C0(n1515), .Y(n947) );
  OAI221X1 U13638 ( .A0(\xArray[3][9] ), .A1(n8284), .B0(\xArray[7][9] ), .B1(
        n8230), .C0(n2241), .Y(n1514) );
  OA22X1 U13639 ( .A0(\xArray[15][9] ), .A1(n8190), .B0(\xArray[11][9] ), .B1(
        n8264), .Y(n2241) );
  OAI221X1 U13640 ( .A0(\xArray[5][8] ), .A1(n8281), .B0(\xArray[9][8] ), .B1(
        n8227), .C0(n1719), .Y(n1252) );
  OAI221X1 U13641 ( .A0(\xArray[5][9] ), .A1(n8281), .B0(\xArray[9][9] ), .B1(
        n8227), .C0(n1716), .Y(n1247) );
  OAI221XL U13642 ( .A0(\xArray[9][7] ), .A1(n8290), .B0(\xArray[13][7] ), 
        .B1(n8236), .C0(n954), .Y(n718) );
  OAI221XL U13643 ( .A0(\xArray[9][8] ), .A1(n8290), .B0(\xArray[13][8] ), 
        .B1(n8236), .C0(n951), .Y(n710) );
  OAI221XL U13644 ( .A0(\xArray[2][5] ), .A1(n8284), .B0(\xArray[6][5] ), .B1(
        n8230), .C0(n2275), .Y(n1727) );
  OAI221XL U13645 ( .A0(\xArray[2][6] ), .A1(n8284), .B0(\xArray[6][6] ), .B1(
        n8230), .C0(n2266), .Y(n1724) );
  OAI221XL U13646 ( .A0(n7463), .A1(n8066), .B0(n7519), .B1(n8063), .C0(n3173), 
        .Y(N28301) );
  OAI221XL U13647 ( .A0(n7463), .A1(n8143), .B0(n7519), .B1(n8140), .C0(n2638), 
        .Y(N28685) );
  OAI221XL U13648 ( .A0(n7465), .A1(n8066), .B0(n7518), .B1(n8063), .C0(n3172), 
        .Y(N28302) );
  OAI221XL U13649 ( .A0(n7465), .A1(n8143), .B0(n7518), .B1(n8140), .C0(n2636), 
        .Y(N28686) );
  OAI221XL U13650 ( .A0(n7467), .A1(n8066), .B0(n7517), .B1(n8063), .C0(n3171), 
        .Y(N28303) );
  OAI221XL U13651 ( .A0(n7467), .A1(n8143), .B0(n7517), .B1(n8140), .C0(n2634), 
        .Y(N28687) );
  OAI221XL U13652 ( .A0(n7469), .A1(n8064), .B0(n7516), .B1(n8063), .C0(n3170), 
        .Y(N28304) );
  OAI221XL U13653 ( .A0(n7469), .A1(n8141), .B0(n7516), .B1(n8140), .C0(n2632), 
        .Y(N28688) );
  OAI221XL U13654 ( .A0(n7471), .A1(n8064), .B0(n7515), .B1(n8063), .C0(n3169), 
        .Y(N28305) );
  OAI221XL U13655 ( .A0(n7471), .A1(n8141), .B0(n7515), .B1(n8140), .C0(n2630), 
        .Y(N28689) );
  OAI22X1 U13656 ( .A0(\xArray[7][44] ), .A1(n7849), .B0(n7861), .B1(n7462), 
        .Y(n3103) );
  OAI22X1 U13657 ( .A0(\xArray[7][45] ), .A1(n7849), .B0(n7861), .B1(n7464), 
        .Y(n3102) );
  OAI22X1 U13658 ( .A0(\xArray[7][46] ), .A1(n7849), .B0(n7862), .B1(n7466), 
        .Y(n3101) );
  OAI22X1 U13659 ( .A0(\xArray[7][47] ), .A1(n7850), .B0(n7862), .B1(n7468), 
        .Y(n3100) );
  OAI22X1 U13660 ( .A0(\xArray[7][48] ), .A1(n7849), .B0(n7862), .B1(n7470), 
        .Y(n3099) );
  OAI22X1 U13661 ( .A0(\xArray[6][44] ), .A1(n7808), .B0(n7821), .B1(n7462), 
        .Y(n3032) );
  OAI22X1 U13662 ( .A0(\xArray[6][45] ), .A1(n7808), .B0(n7822), .B1(n7464), 
        .Y(n3031) );
  OAI22X1 U13663 ( .A0(\xArray[6][46] ), .A1(n7808), .B0(n7820), .B1(n7466), 
        .Y(n3030) );
  OAI22X1 U13664 ( .A0(\xArray[6][47] ), .A1(n7808), .B0(n7822), .B1(n7468), 
        .Y(n3029) );
  OAI22X1 U13665 ( .A0(\xArray[6][48] ), .A1(n7808), .B0(n7821), .B1(n7470), 
        .Y(n3028) );
  AND4X1 U13666 ( .A(n4029), .B(n4030), .C(n4031), .D(n4032), .Y(n2388) );
  AOI221XL U13667 ( .A0(n7964), .A1(\xArray[9][44] ), .B0(\xArray[8][44] ), 
        .B1(n7960), .C0(n4033), .Y(n4032) );
  AOI221XL U13668 ( .A0(n7948), .A1(n7462), .B0(n7945), .B1(\xArray[2][44] ), 
        .C0(n4035), .Y(n4031) );
  AND4X1 U13669 ( .A(n4011), .B(n4012), .C(n4013), .D(n4014), .Y(n2385) );
  AOI221XL U13670 ( .A0(n7964), .A1(\xArray[9][45] ), .B0(\xArray[8][45] ), 
        .B1(n7960), .C0(n4015), .Y(n4014) );
  AOI221XL U13671 ( .A0(n7948), .A1(n7464), .B0(n7945), .B1(\xArray[2][45] ), 
        .C0(n4017), .Y(n4013) );
  AND4X1 U13672 ( .A(n3993), .B(n3994), .C(n3995), .D(n3996), .Y(n2382) );
  AOI221XL U13673 ( .A0(n7964), .A1(\xArray[9][46] ), .B0(\xArray[8][46] ), 
        .B1(n7960), .C0(n3997), .Y(n3996) );
  AOI221XL U13674 ( .A0(n7948), .A1(n7466), .B0(n7945), .B1(\xArray[2][46] ), 
        .C0(n3999), .Y(n3995) );
  AND4X1 U13675 ( .A(n3975), .B(n3976), .C(n3977), .D(n3978), .Y(n2379) );
  AOI221XL U13676 ( .A0(n7964), .A1(\xArray[9][47] ), .B0(\xArray[8][47] ), 
        .B1(n7960), .C0(n3979), .Y(n3978) );
  AOI221XL U13677 ( .A0(n7948), .A1(n7468), .B0(n7945), .B1(\xArray[2][47] ), 
        .C0(n3981), .Y(n3977) );
  AND4X1 U13678 ( .A(n3957), .B(n3958), .C(n3959), .D(n3960), .Y(n2376) );
  AOI221XL U13679 ( .A0(n7964), .A1(\xArray[9][48] ), .B0(\xArray[8][48] ), 
        .B1(n7960), .C0(n3961), .Y(n3960) );
  AOI221XL U13680 ( .A0(n7948), .A1(n7470), .B0(n7945), .B1(\xArray[2][48] ), 
        .C0(n3963), .Y(n3959) );
  AOI221XL U13681 ( .A0(\xArray[13][1] ), .A1(n1746), .B0(\xArray[1][1] ), 
        .B1(n1747), .C0(n2308), .Y(n2307) );
  OA22X1 U13682 ( .A0(n8323), .A1(n1546), .B0(n7728), .B1(n1739), .Y(n2306) );
  OAI22XL U13683 ( .A0(n8175), .A1(n9388), .B0(n8171), .B1(n9386), .Y(n2308)
         );
  AOI221XL U13684 ( .A0(\xArray[13][2] ), .A1(n8180), .B0(\xArray[1][2] ), 
        .B1(n8176), .C0(n2299), .Y(n2298) );
  OAI22XL U13685 ( .A0(n8175), .A1(n9380), .B0(n8171), .B1(n9378), .Y(n2299)
         );
  AOI221XL U13686 ( .A0(\xArray[13][3] ), .A1(n8180), .B0(\xArray[1][3] ), 
        .B1(n8176), .C0(n2290), .Y(n2289) );
  OAI22XL U13687 ( .A0(n8175), .A1(n9372), .B0(n8171), .B1(n9370), .Y(n2290)
         );
  OAI221X1 U13688 ( .A0(\xArray[7][10] ), .A1(n8296), .B0(\xArray[11][10] ), 
        .B1(n8242), .C0(n1244), .Y(n693) );
  OAI221X1 U13689 ( .A0(\xArray[7][11] ), .A1(n8296), .B0(\xArray[11][11] ), 
        .B1(n8242), .C0(n1239), .Y(n685) );
  AOI2BB2X1 U13690 ( .B0(n9304), .B1(n8212), .A0N(\xArray[15][11] ), .A1N(
        n8255), .Y(n1239) );
  OAI221X1 U13691 ( .A0(\xArray[4][10] ), .A1(n8284), .B0(\xArray[8][10] ), 
        .B1(n8230), .C0(n2233), .Y(n1508) );
  OA22X1 U13692 ( .A0(\xArray[0][10] ), .A1(n8190), .B0(\xArray[12][10] ), 
        .B1(n8264), .Y(n2233) );
  OAI221X1 U13693 ( .A0(\xArray[4][11] ), .A1(n8285), .B0(\xArray[8][11] ), 
        .B1(n8231), .C0(n2224), .Y(n1504) );
  OA22X1 U13694 ( .A0(\xArray[0][11] ), .A1(n8190), .B0(\xArray[12][11] ), 
        .B1(n8264), .Y(n2224) );
  OAI221X1 U13695 ( .A0(\xArray[8][9] ), .A1(n8296), .B0(\xArray[12][9] ), 
        .B1(n8242), .C0(n1248), .Y(n703) );
  OAI221X1 U13696 ( .A0(\xArray[8][10] ), .A1(n8296), .B0(\xArray[12][10] ), 
        .B1(n8242), .C0(n1243), .Y(n695) );
  OAI221X1 U13697 ( .A0(\xArray[6][10] ), .A1(n8293), .B0(\xArray[10][10] ), 
        .B1(n8239), .C0(n1511), .Y(n944) );
  OA22X1 U13698 ( .A0(\xArray[14][10] ), .A1(n8272), .B0(\xArray[2][10] ), 
        .B1(n8186), .Y(n1511) );
  OAI221X1 U13699 ( .A0(\xArray[3][10] ), .A1(n8284), .B0(\xArray[7][10] ), 
        .B1(n8230), .C0(n2232), .Y(n1510) );
  OA22X1 U13700 ( .A0(\xArray[15][10] ), .A1(n8190), .B0(\xArray[11][10] ), 
        .B1(n8264), .Y(n2232) );
  OAI221X1 U13701 ( .A0(\xArray[6][11] ), .A1(n8293), .B0(\xArray[10][11] ), 
        .B1(n8239), .C0(n1507), .Y(n941) );
  OAI221X1 U13702 ( .A0(\xArray[3][11] ), .A1(n8285), .B0(\xArray[7][11] ), 
        .B1(n8231), .C0(n2223), .Y(n1506) );
  OA22X1 U13703 ( .A0(\xArray[15][11] ), .A1(n8190), .B0(\xArray[11][11] ), 
        .B1(n8264), .Y(n2223) );
  OAI221X1 U13704 ( .A0(\xArray[5][10] ), .A1(n8281), .B0(\xArray[9][10] ), 
        .B1(n8227), .C0(n1713), .Y(n1242) );
  OAI221X1 U13705 ( .A0(\xArray[5][11] ), .A1(n8281), .B0(\xArray[9][11] ), 
        .B1(n8227), .C0(n1710), .Y(n1237) );
  OAI221XL U13706 ( .A0(\xArray[9][9] ), .A1(n8290), .B0(\xArray[13][9] ), 
        .B1(n8236), .C0(n948), .Y(n702) );
  OAI221XL U13707 ( .A0(\xArray[9][10] ), .A1(n8290), .B0(\xArray[13][10] ), 
        .B1(n8236), .C0(n945), .Y(n694) );
  OAI221XL U13708 ( .A0(\xArray[2][7] ), .A1(n8284), .B0(\xArray[6][7] ), .B1(
        n8230), .C0(n2257), .Y(n1721) );
  OAI221XL U13709 ( .A0(\xArray[2][8] ), .A1(n8284), .B0(\xArray[6][8] ), .B1(
        n8230), .C0(n2248), .Y(n1718) );
  AOI221XL U13710 ( .A0(n7948), .A1(n7457), .B0(n7945), .B1(\xArray[2][41] ), 
        .C0(n4089), .Y(n4085) );
  OAI222XL U13711 ( .A0(n9066), .A1(n7942), .B0(n8558), .B1(n7939), .C0(n7936), 
        .C1(n9065), .Y(n4089) );
  AOI221XL U13712 ( .A0(n7948), .A1(n7459), .B0(n7945), .B1(\xArray[2][42] ), 
        .C0(n4071), .Y(n4067) );
  OAI222XL U13713 ( .A0(n9058), .A1(n7942), .B0(n8553), .B1(n7939), .C0(n7936), 
        .C1(n9057), .Y(n4071) );
  OAI221XL U13714 ( .A0(n7458), .A1(n8064), .B0(n7522), .B1(n8063), .C0(n3176), 
        .Y(N28298) );
  OAI221XL U13715 ( .A0(n7458), .A1(n8141), .B0(n7522), .B1(n8140), .C0(n2644), 
        .Y(N28682) );
  OAI221XL U13716 ( .A0(n7460), .A1(n6607), .B0(n7521), .B1(n8063), .C0(n3175), 
        .Y(N28299) );
  OAI221XL U13717 ( .A0(n7460), .A1(n6608), .B0(n7521), .B1(n8140), .C0(n2642), 
        .Y(N28683) );
  OAI221XL U13718 ( .A0(n6623), .A1(n6607), .B0(n7520), .B1(n8063), .C0(n3174), 
        .Y(N28300) );
  OAI221XL U13719 ( .A0(n6623), .A1(n6608), .B0(n7520), .B1(n8140), .C0(n2640), 
        .Y(N28684) );
  AOI221XL U13720 ( .A0(n7964), .A1(\xArray[9][43] ), .B0(\xArray[8][43] ), 
        .B1(n7960), .C0(n4051), .Y(n4050) );
  AOI221XL U13721 ( .A0(n7948), .A1(n7461), .B0(n7945), .B1(\xArray[2][43] ), 
        .C0(n4053), .Y(n4049) );
  AOI221XL U13722 ( .A0(\xArray[13][0] ), .A1(n1746), .B0(\xArray[1][0] ), 
        .B1(n1747), .C0(n2317), .Y(n2316) );
  OAI22XL U13723 ( .A0(n8175), .A1(n9396), .B0(n8171), .B1(n9394), .Y(n2317)
         );
  OAI221X1 U13724 ( .A0(\xArray[7][12] ), .A1(n8296), .B0(\xArray[11][12] ), 
        .B1(n8242), .C0(n1234), .Y(n677) );
  AOI2BB2X1 U13725 ( .B0(n9296), .B1(n8212), .A0N(\xArray[15][12] ), .A1N(
        n8255), .Y(n1234) );
  OAI221X1 U13726 ( .A0(\xArray[7][13] ), .A1(n8296), .B0(\xArray[11][13] ), 
        .B1(n8242), .C0(n1229), .Y(n669) );
  AOI2BB2X1 U13727 ( .B0(n9288), .B1(n8212), .A0N(\xArray[15][13] ), .A1N(
        n8255), .Y(n1229) );
  OAI221X1 U13728 ( .A0(\xArray[4][12] ), .A1(n8285), .B0(\xArray[8][12] ), 
        .B1(n8231), .C0(n2215), .Y(n1500) );
  OAI221X1 U13729 ( .A0(\xArray[4][13] ), .A1(n8285), .B0(\xArray[8][13] ), 
        .B1(n8231), .C0(n2206), .Y(n1496) );
  OAI221X1 U13730 ( .A0(\xArray[8][11] ), .A1(n8296), .B0(\xArray[12][11] ), 
        .B1(n8242), .C0(n1238), .Y(n687) );
  OAI221X1 U13731 ( .A0(\xArray[8][12] ), .A1(n8296), .B0(\xArray[12][12] ), 
        .B1(n8242), .C0(n1233), .Y(n679) );
  OAI221X1 U13732 ( .A0(\xArray[6][12] ), .A1(n8293), .B0(\xArray[10][12] ), 
        .B1(n8239), .C0(n1503), .Y(n938) );
  OAI221X1 U13733 ( .A0(\xArray[3][12] ), .A1(n8285), .B0(\xArray[7][12] ), 
        .B1(n8231), .C0(n2214), .Y(n1502) );
  OAI221X1 U13734 ( .A0(\xArray[6][13] ), .A1(n8293), .B0(\xArray[10][13] ), 
        .B1(n8239), .C0(n1499), .Y(n935) );
  OAI221X1 U13735 ( .A0(\xArray[3][13] ), .A1(n8285), .B0(\xArray[7][13] ), 
        .B1(n8231), .C0(n2205), .Y(n1498) );
  OAI221X1 U13736 ( .A0(\xArray[5][12] ), .A1(n8281), .B0(\xArray[9][12] ), 
        .B1(n8227), .C0(n1707), .Y(n1232) );
  OAI221X1 U13737 ( .A0(\xArray[5][13] ), .A1(n8281), .B0(\xArray[9][13] ), 
        .B1(n8227), .C0(n1704), .Y(n1227) );
  OAI221XL U13738 ( .A0(\xArray[9][11] ), .A1(n8290), .B0(\xArray[13][11] ), 
        .B1(n8236), .C0(n942), .Y(n686) );
  OAI221XL U13739 ( .A0(\xArray[9][12] ), .A1(n8290), .B0(\xArray[13][12] ), 
        .B1(n8236), .C0(n939), .Y(n678) );
  OAI221XL U13740 ( .A0(\xArray[2][9] ), .A1(n8284), .B0(\xArray[6][9] ), .B1(
        n8230), .C0(n2239), .Y(n1715) );
  OAI221XL U13741 ( .A0(\xArray[2][10] ), .A1(n8284), .B0(\xArray[6][10] ), 
        .B1(n8230), .C0(n2230), .Y(n1712) );
  OAI221XL U13742 ( .A0(n7448), .A1(n8066), .B0(n7527), .B1(n8063), .C0(n3181), 
        .Y(N28293) );
  OAI221XL U13743 ( .A0(n7448), .A1(n8143), .B0(n7527), .B1(n8138), .C0(n2654), 
        .Y(N28677) );
  OAI221XL U13744 ( .A0(n7450), .A1(n8066), .B0(n7526), .B1(n8063), .C0(n3180), 
        .Y(N28294) );
  OAI221XL U13745 ( .A0(n7450), .A1(n8143), .B0(n7526), .B1(n8138), .C0(n2652), 
        .Y(N28678) );
  OAI221XL U13746 ( .A0(n7452), .A1(n8066), .B0(n7525), .B1(n8063), .C0(n3179), 
        .Y(N28295) );
  OAI221XL U13747 ( .A0(n7452), .A1(n8143), .B0(n7525), .B1(n8140), .C0(n2650), 
        .Y(N28679) );
  OAI221XL U13748 ( .A0(n7454), .A1(n8066), .B0(n7524), .B1(n8063), .C0(n3178), 
        .Y(N28296) );
  OAI221XL U13749 ( .A0(n7454), .A1(n8143), .B0(n7524), .B1(n8140), .C0(n2648), 
        .Y(N28680) );
  OAI221XL U13750 ( .A0(n7456), .A1(n6607), .B0(n7523), .B1(n8063), .C0(n3177), 
        .Y(N28297) );
  OAI221XL U13751 ( .A0(n7456), .A1(n6608), .B0(n7523), .B1(n8140), .C0(n2646), 
        .Y(N28681) );
  OAI22X1 U13752 ( .A0(\xArray[7][36] ), .A1(n7848), .B0(n7863), .B1(n7447), 
        .Y(n3111) );
  OAI22X1 U13753 ( .A0(\xArray[7][37] ), .A1(n7848), .B0(n7864), .B1(n7449), 
        .Y(n3110) );
  OAI22X1 U13754 ( .A0(\xArray[7][38] ), .A1(n7848), .B0(n7860), .B1(n7451), 
        .Y(n3109) );
  OAI22X1 U13755 ( .A0(\xArray[7][39] ), .A1(n7848), .B0(n7860), .B1(n7453), 
        .Y(n3108) );
  OAI22X1 U13756 ( .A0(\xArray[7][40] ), .A1(n7849), .B0(n7860), .B1(n7455), 
        .Y(n3107) );
  OAI22X1 U13757 ( .A0(\xArray[6][36] ), .A1(n7809), .B0(n7820), .B1(n7447), 
        .Y(n3040) );
  OAI22X1 U13758 ( .A0(\xArray[6][37] ), .A1(n7809), .B0(n7820), .B1(n7449), 
        .Y(n3039) );
  OAI22X1 U13759 ( .A0(\xArray[6][38] ), .A1(n7809), .B0(n7822), .B1(n7451), 
        .Y(n3038) );
  OAI22X1 U13760 ( .A0(\xArray[6][39] ), .A1(n7809), .B0(n7822), .B1(n7453), 
        .Y(n3037) );
  OAI22X1 U13761 ( .A0(\xArray[6][40] ), .A1(n7808), .B0(n7821), .B1(n7455), 
        .Y(n3036) );
  AND4X1 U13762 ( .A(n4173), .B(n4174), .C(n4175), .D(n4176), .Y(n2412) );
  AOI221XL U13763 ( .A0(n7965), .A1(\xArray[9][36] ), .B0(\xArray[8][36] ), 
        .B1(n7961), .C0(n4177), .Y(n4176) );
  AOI221XL U13764 ( .A0(n7947), .A1(n7447), .B0(n7944), .B1(\xArray[2][36] ), 
        .C0(n4179), .Y(n4175) );
  AND4X1 U13765 ( .A(n4155), .B(n4156), .C(n4157), .D(n4158), .Y(n2409) );
  AOI221XL U13766 ( .A0(n7965), .A1(\xArray[9][37] ), .B0(\xArray[8][37] ), 
        .B1(n7961), .C0(n4159), .Y(n4158) );
  AOI221XL U13767 ( .A0(n7948), .A1(n7449), .B0(n7944), .B1(\xArray[2][37] ), 
        .C0(n4161), .Y(n4157) );
  AND4X1 U13768 ( .A(n4137), .B(n4138), .C(n4139), .D(n4140), .Y(n2406) );
  AOI221XL U13769 ( .A0(n7965), .A1(\xArray[9][38] ), .B0(\xArray[8][38] ), 
        .B1(n7961), .C0(n4141), .Y(n4140) );
  AOI221XL U13770 ( .A0(n7949), .A1(n7451), .B0(n7944), .B1(\xArray[2][38] ), 
        .C0(n4143), .Y(n4139) );
  AND4X1 U13771 ( .A(n4119), .B(n4120), .C(n4121), .D(n4122), .Y(n2403) );
  AOI221XL U13772 ( .A0(n7965), .A1(\xArray[9][39] ), .B0(\xArray[8][39] ), 
        .B1(n7961), .C0(n4123), .Y(n4122) );
  AOI221XL U13773 ( .A0(n7947), .A1(n7453), .B0(n7944), .B1(\xArray[2][39] ), 
        .C0(n4125), .Y(n4121) );
  AND4X1 U13774 ( .A(n4101), .B(n4102), .C(n4103), .D(n4104), .Y(n2400) );
  AOI221XL U13775 ( .A0(n7964), .A1(\xArray[9][40] ), .B0(\xArray[8][40] ), 
        .B1(n7960), .C0(n4105), .Y(n4104) );
  AOI221XL U13776 ( .A0(n7948), .A1(n7455), .B0(n7945), .B1(\xArray[2][40] ), 
        .C0(n4107), .Y(n4103) );
  AOI221XL U13777 ( .A0(\xArray[13][4] ), .A1(n8180), .B0(\xArray[1][4] ), 
        .B1(n8178), .C0(n2281), .Y(n2280) );
  OAI22XL U13778 ( .A0(n8175), .A1(n9364), .B0(n8171), .B1(n9362), .Y(n2281)
         );
  AOI221XL U13779 ( .A0(\xArray[13][5] ), .A1(n8180), .B0(\xArray[1][5] ), 
        .B1(n8178), .C0(n2272), .Y(n2271) );
  OAI22XL U13780 ( .A0(n8175), .A1(n9356), .B0(n8171), .B1(n9354), .Y(n2272)
         );
  AOI221XL U13781 ( .A0(\xArray[13][6] ), .A1(n8180), .B0(\xArray[1][6] ), 
        .B1(n8178), .C0(n2263), .Y(n2262) );
  OAI22XL U13782 ( .A0(n8175), .A1(n9348), .B0(n8171), .B1(n9346), .Y(n2263)
         );
  AOI221XL U13783 ( .A0(\xArray[13][7] ), .A1(n1746), .B0(\xArray[1][7] ), 
        .B1(n8178), .C0(n2254), .Y(n2253) );
  OAI22XL U13784 ( .A0(n8175), .A1(n9340), .B0(n8171), .B1(n9338), .Y(n2254)
         );
  OAI221X1 U13785 ( .A0(\xArray[7][14] ), .A1(n8296), .B0(\xArray[11][14] ), 
        .B1(n8242), .C0(n1224), .Y(n661) );
  AOI2BB2X1 U13786 ( .B0(n9280), .B1(n8212), .A0N(\xArray[15][14] ), .A1N(
        n8255), .Y(n1224) );
  OAI221X1 U13787 ( .A0(\xArray[4][14] ), .A1(n8285), .B0(\xArray[8][14] ), 
        .B1(n8231), .C0(n2197), .Y(n1492) );
  OAI221X1 U13788 ( .A0(\xArray[4][15] ), .A1(n8285), .B0(\xArray[8][15] ), 
        .B1(n8231), .C0(n2188), .Y(n1488) );
  OAI221X1 U13789 ( .A0(\xArray[8][13] ), .A1(n8296), .B0(\xArray[12][13] ), 
        .B1(n8242), .C0(n1228), .Y(n671) );
  OAI221X1 U13790 ( .A0(\xArray[8][14] ), .A1(n8296), .B0(\xArray[12][14] ), 
        .B1(n8242), .C0(n1223), .Y(n663) );
  OAI221X1 U13791 ( .A0(\xArray[6][14] ), .A1(n8293), .B0(\xArray[10][14] ), 
        .B1(n8239), .C0(n1495), .Y(n932) );
  OAI221X1 U13792 ( .A0(\xArray[3][14] ), .A1(n8285), .B0(\xArray[7][14] ), 
        .B1(n8231), .C0(n2196), .Y(n1494) );
  OAI221X1 U13793 ( .A0(\xArray[6][15] ), .A1(n8293), .B0(\xArray[10][15] ), 
        .B1(n8239), .C0(n1491), .Y(n929) );
  OAI221X1 U13794 ( .A0(\xArray[3][15] ), .A1(n8285), .B0(\xArray[7][15] ), 
        .B1(n8231), .C0(n2187), .Y(n1490) );
  OAI221X1 U13795 ( .A0(\xArray[5][14] ), .A1(n8281), .B0(\xArray[9][14] ), 
        .B1(n8227), .C0(n1701), .Y(n1222) );
  OA22X1 U13796 ( .A0(\xArray[1][14] ), .A1(n8188), .B0(\xArray[13][14] ), 
        .B1(n8259), .Y(n1701) );
  OAI221X1 U13797 ( .A0(\xArray[5][15] ), .A1(n8281), .B0(\xArray[9][15] ), 
        .B1(n8227), .C0(n1698), .Y(n1217) );
  OA22X1 U13798 ( .A0(\xArray[1][15] ), .A1(n8188), .B0(\xArray[13][15] ), 
        .B1(n8259), .Y(n1698) );
  NAND2BX2 U13799 ( .AN(n768), .B(n769), .Y(N34026) );
  OAI222XL U13800 ( .A0(n780), .A1(n8340), .B0(n781), .B1(n8308), .C0(n782), 
        .C1(n7712), .Y(n768) );
  AOI221XL U13801 ( .A0(\xArray[14][0] ), .A1(n6573), .B0(\xArray[2][0] ), 
        .B1(n8362), .C0(n770), .Y(n769) );
  OAI22XL U13802 ( .A0(n8357), .A1(n9395), .B0(n8355), .B1(n9397), .Y(n770) );
  OAI221XL U13803 ( .A0(\xArray[9][13] ), .A1(n8290), .B0(\xArray[13][13] ), 
        .B1(n8236), .C0(n936), .Y(n670) );
  OAI221XL U13804 ( .A0(\xArray[9][14] ), .A1(n8290), .B0(\xArray[13][14] ), 
        .B1(n8236), .C0(n933), .Y(n662) );
  OAI221XL U13805 ( .A0(\xArray[2][11] ), .A1(n8285), .B0(\xArray[6][11] ), 
        .B1(n8231), .C0(n2221), .Y(n1709) );
  OAI221XL U13806 ( .A0(\xArray[2][12] ), .A1(n8285), .B0(\xArray[6][12] ), 
        .B1(n8231), .C0(n2212), .Y(n1706) );
  NAND2BX2 U13807 ( .AN(n760), .B(n761), .Y(N34027) );
  OAI222XL U13808 ( .A0(n765), .A1(n8340), .B0(n766), .B1(n8308), .C0(n767), 
        .C1(n7712), .Y(n760) );
  AOI221XL U13809 ( .A0(\xArray[14][1] ), .A1(n6573), .B0(\xArray[2][1] ), 
        .B1(n8362), .C0(n762), .Y(n761) );
  OAI22XL U13810 ( .A0(n8357), .A1(n9387), .B0(n8355), .B1(n9389), .Y(n762) );
  OAI222XL U13811 ( .A0(n757), .A1(n8340), .B0(n758), .B1(n8308), .C0(n759), 
        .C1(n7712), .Y(n752) );
  AOI221XL U13812 ( .A0(\xArray[14][2] ), .A1(n6573), .B0(\xArray[2][2] ), 
        .B1(n8362), .C0(n754), .Y(n753) );
  OAI22XL U13813 ( .A0(n8357), .A1(n9379), .B0(n8355), .B1(n9381), .Y(n754) );
  OAI222XL U13814 ( .A0(n749), .A1(n8340), .B0(n750), .B1(n8308), .C0(n751), 
        .C1(n7712), .Y(n744) );
  AOI221XL U13815 ( .A0(\xArray[14][3] ), .A1(n6573), .B0(\xArray[2][3] ), 
        .B1(n8362), .C0(n746), .Y(n745) );
  OAI22XL U13816 ( .A0(n8357), .A1(n9371), .B0(n8355), .B1(n9373), .Y(n746) );
  AOI221XL U13817 ( .A0(n7948), .A1(n7439), .B0(n7944), .B1(\xArray[2][32] ), 
        .C0(n4251), .Y(n4247) );
  OAI222XL U13818 ( .A0(n9138), .A1(n7943), .B0(n8603), .B1(n7940), .C0(n7937), 
        .C1(n9137), .Y(n4251) );
  OAI221XL U13819 ( .A0(n7440), .A1(n8066), .B0(n7531), .B1(n8061), .C0(n3185), 
        .Y(N28289) );
  OAI221XL U13820 ( .A0(n7440), .A1(n8143), .B0(n7531), .B1(n8139), .C0(n2662), 
        .Y(N28673) );
  OAI221XL U13821 ( .A0(n7442), .A1(n8066), .B0(n7530), .B1(n8061), .C0(n3184), 
        .Y(N28290) );
  OAI221XL U13822 ( .A0(n7442), .A1(n8143), .B0(n7530), .B1(n8139), .C0(n2660), 
        .Y(N28674) );
  OAI221XL U13823 ( .A0(n7444), .A1(n8066), .B0(n7529), .B1(n8061), .C0(n3183), 
        .Y(N28291) );
  OAI221XL U13824 ( .A0(n7444), .A1(n8143), .B0(n7529), .B1(n8140), .C0(n2658), 
        .Y(N28675) );
  OAI221XL U13825 ( .A0(n7446), .A1(n8066), .B0(n7528), .B1(n8061), .C0(n3182), 
        .Y(N28292) );
  OAI221XL U13826 ( .A0(n7446), .A1(n8143), .B0(n7528), .B1(n8140), .C0(n2656), 
        .Y(N28676) );
  OAI22X1 U13827 ( .A0(\xArray[7][33] ), .A1(n7848), .B0(n7859), .B1(n7441), 
        .Y(n3114) );
  OAI22X1 U13828 ( .A0(\xArray[7][34] ), .A1(n7848), .B0(n7864), .B1(n7443), 
        .Y(n3113) );
  OAI22X1 U13829 ( .A0(\xArray[7][35] ), .A1(n7848), .B0(n7863), .B1(n7445), 
        .Y(n3112) );
  OAI22X1 U13830 ( .A0(\xArray[6][33] ), .A1(n7809), .B0(n7819), .B1(n7441), 
        .Y(n3043) );
  OAI22X1 U13831 ( .A0(\xArray[6][34] ), .A1(n7809), .B0(n7820), .B1(n7443), 
        .Y(n3042) );
  OAI22X1 U13832 ( .A0(\xArray[6][35] ), .A1(n7809), .B0(n7820), .B1(n7445), 
        .Y(n3041) );
  AND4X1 U13833 ( .A(n4227), .B(n4228), .C(n4229), .D(n4230), .Y(n2421) );
  AOI221XL U13834 ( .A0(n7965), .A1(\xArray[9][33] ), .B0(\xArray[8][33] ), 
        .B1(n7961), .C0(n4231), .Y(n4230) );
  AOI221XL U13835 ( .A0(n7948), .A1(n7441), .B0(n7944), .B1(\xArray[2][33] ), 
        .C0(n4233), .Y(n4229) );
  AND4X1 U13836 ( .A(n4209), .B(n4210), .C(n4211), .D(n4212), .Y(n2418) );
  AOI221XL U13837 ( .A0(n7965), .A1(\xArray[9][34] ), .B0(\xArray[8][34] ), 
        .B1(n7961), .C0(n4213), .Y(n4212) );
  AOI221XL U13838 ( .A0(n7949), .A1(n7443), .B0(n7944), .B1(\xArray[2][34] ), 
        .C0(n4215), .Y(n4211) );
  AND4X1 U13839 ( .A(n4191), .B(n4192), .C(n4193), .D(n4194), .Y(n2415) );
  AOI221XL U13840 ( .A0(n7965), .A1(\xArray[9][35] ), .B0(\xArray[8][35] ), 
        .B1(n7961), .C0(n4195), .Y(n4194) );
  AOI221XL U13841 ( .A0(n7947), .A1(n7445), .B0(n3667), .B1(\xArray[2][35] ), 
        .C0(n4197), .Y(n4193) );
  OAI221X1 U13842 ( .A0(\xArray[7][15] ), .A1(n8296), .B0(\xArray[11][15] ), 
        .B1(n8242), .C0(n1219), .Y(n653) );
  AOI2BB2X1 U13843 ( .B0(n9272), .B1(n8212), .A0N(\xArray[15][15] ), .A1N(
        n8255), .Y(n1219) );
  OAI221X1 U13844 ( .A0(\xArray[7][16] ), .A1(n8296), .B0(\xArray[11][16] ), 
        .B1(n8242), .C0(n1214), .Y(n645) );
  AOI2BB2X1 U13845 ( .B0(n9264), .B1(n8212), .A0N(\xArray[15][16] ), .A1N(
        n8255), .Y(n1214) );
  OAI221X1 U13846 ( .A0(\xArray[4][17] ), .A1(n8286), .B0(\xArray[8][17] ), 
        .B1(n8232), .C0(n2170), .Y(n1480) );
  OA22X1 U13847 ( .A0(\xArray[0][17] ), .A1(n8191), .B0(\xArray[12][17] ), 
        .B1(n8265), .Y(n2170) );
  OAI221X1 U13848 ( .A0(\xArray[8][15] ), .A1(n8296), .B0(\xArray[12][15] ), 
        .B1(n8242), .C0(n1218), .Y(n655) );
  OAI221X1 U13849 ( .A0(\xArray[8][16] ), .A1(n8296), .B0(\xArray[12][16] ), 
        .B1(n8242), .C0(n1213), .Y(n647) );
  OAI221X1 U13850 ( .A0(\xArray[6][16] ), .A1(n8293), .B0(\xArray[10][16] ), 
        .B1(n8239), .C0(n1487), .Y(n926) );
  OAI221X1 U13851 ( .A0(\xArray[3][16] ), .A1(n8285), .B0(\xArray[7][16] ), 
        .B1(n8231), .C0(n2178), .Y(n1486) );
  OA22X1 U13852 ( .A0(\xArray[15][16] ), .A1(n8191), .B0(\xArray[11][16] ), 
        .B1(n8265), .Y(n2178) );
  OAI221X1 U13853 ( .A0(\xArray[3][17] ), .A1(n8286), .B0(\xArray[7][17] ), 
        .B1(n8232), .C0(n2169), .Y(n1482) );
  OA22X1 U13854 ( .A0(\xArray[15][17] ), .A1(n8191), .B0(\xArray[11][17] ), 
        .B1(n8265), .Y(n2169) );
  OAI221X1 U13855 ( .A0(\xArray[5][16] ), .A1(n8281), .B0(\xArray[9][16] ), 
        .B1(n8227), .C0(n1695), .Y(n1212) );
  OA22X1 U13856 ( .A0(\xArray[1][16] ), .A1(n8188), .B0(\xArray[13][16] ), 
        .B1(n8259), .Y(n1695) );
  OAI221X1 U13857 ( .A0(\xArray[5][17] ), .A1(n8281), .B0(\xArray[9][17] ), 
        .B1(n8227), .C0(n1692), .Y(n1207) );
  OAI221XL U13858 ( .A0(\xArray[9][15] ), .A1(n8290), .B0(\xArray[13][15] ), 
        .B1(n8236), .C0(n930), .Y(n654) );
  OAI221XL U13859 ( .A0(\xArray[9][16] ), .A1(n8290), .B0(\xArray[13][16] ), 
        .B1(n8236), .C0(n927), .Y(n646) );
  OA22X1 U13860 ( .A0(\xArray[5][16] ), .A1(n8195), .B0(\xArray[1][16] ), .B1(
        n8269), .Y(n927) );
  OAI221XL U13861 ( .A0(\xArray[2][14] ), .A1(n8285), .B0(\xArray[6][14] ), 
        .B1(n8231), .C0(n2194), .Y(n1700) );
  AOI221XL U13862 ( .A0(n7947), .A1(n7437), .B0(n7944), .B1(\xArray[2][31] ), 
        .C0(n4269), .Y(n4265) );
  OAI222XL U13863 ( .A0(n9146), .A1(n7943), .B0(n8608), .B1(n7940), .C0(n7937), 
        .C1(n9145), .Y(n4269) );
  OAI221XL U13864 ( .A0(n7434), .A1(n8066), .B0(n7534), .B1(n8061), .C0(n3188), 
        .Y(N28286) );
  OAI221XL U13865 ( .A0(n7434), .A1(n8143), .B0(n7534), .B1(n8140), .C0(n2668), 
        .Y(N28670) );
  OAI221XL U13866 ( .A0(n7436), .A1(n8066), .B0(n7533), .B1(n8062), .C0(n3187), 
        .Y(N28287) );
  OAI221XL U13867 ( .A0(n7436), .A1(n8143), .B0(n7533), .B1(n8138), .C0(n2666), 
        .Y(N28671) );
  OAI221XL U13868 ( .A0(n7438), .A1(n8066), .B0(n7532), .B1(n8063), .C0(n3186), 
        .Y(N28288) );
  OAI221XL U13869 ( .A0(n7438), .A1(n8143), .B0(n7532), .B1(n8140), .C0(n2664), 
        .Y(N28672) );
  OAI22X1 U13870 ( .A0(\xArray[7][28] ), .A1(n7848), .B0(n7860), .B1(n7431), 
        .Y(n3119) );
  OAI22X1 U13871 ( .A0(\xArray[7][29] ), .A1(n7848), .B0(n7863), .B1(n7433), 
        .Y(n3118) );
  OAI22X1 U13872 ( .A0(\xArray[7][30] ), .A1(n7848), .B0(n7864), .B1(n7435), 
        .Y(n3117) );
  OAI22X1 U13873 ( .A0(\xArray[6][28] ), .A1(n7809), .B0(n7820), .B1(n7431), 
        .Y(n3048) );
  OAI22X1 U13874 ( .A0(\xArray[6][29] ), .A1(n7809), .B0(n7822), .B1(n7433), 
        .Y(n3047) );
  OAI22X1 U13875 ( .A0(\xArray[6][30] ), .A1(n7809), .B0(n7822), .B1(n7435), 
        .Y(n3046) );
  OAI221XL U13876 ( .A0(\xArray[2][13] ), .A1(n8285), .B0(\xArray[6][13] ), 
        .B1(n8231), .C0(n2203), .Y(n1703) );
  CLKBUFX3 U13877 ( .A(n2436), .Y(n7432) );
  AND4X1 U13878 ( .A(n4317), .B(n4318), .C(n4319), .D(n4320), .Y(n2436) );
  AOI221XL U13879 ( .A0(n7965), .A1(\xArray[9][28] ), .B0(\xArray[8][28] ), 
        .B1(n7961), .C0(n4321), .Y(n4320) );
  AOI221XL U13880 ( .A0(n6603), .A1(n7431), .B0(n7944), .B1(\xArray[2][28] ), 
        .C0(n4323), .Y(n4319) );
  AND4X1 U13881 ( .A(n4299), .B(n4300), .C(n4301), .D(n4302), .Y(n2433) );
  AOI221XL U13882 ( .A0(n7965), .A1(\xArray[9][29] ), .B0(\xArray[8][29] ), 
        .B1(n7961), .C0(n4303), .Y(n4302) );
  AOI221XL U13883 ( .A0(n7948), .A1(n7433), .B0(n7945), .B1(\xArray[2][29] ), 
        .C0(n4305), .Y(n4301) );
  AND4X1 U13884 ( .A(n4281), .B(n4282), .C(n4283), .D(n4284), .Y(n2430) );
  AOI221XL U13885 ( .A0(n7965), .A1(\xArray[9][30] ), .B0(\xArray[8][30] ), 
        .B1(n7961), .C0(n4285), .Y(n4284) );
  AOI221XL U13886 ( .A0(n7949), .A1(n7435), .B0(n7946), .B1(\xArray[2][30] ), 
        .C0(n4287), .Y(n4283) );
  AOI221XL U13887 ( .A0(\xArray[13][8] ), .A1(n8180), .B0(\xArray[1][8] ), 
        .B1(n8178), .C0(n2245), .Y(n2244) );
  OAI22XL U13888 ( .A0(n8175), .A1(n9332), .B0(n8171), .B1(n9330), .Y(n2245)
         );
  AOI221XL U13889 ( .A0(\xArray[13][9] ), .A1(n8180), .B0(\xArray[1][9] ), 
        .B1(n8178), .C0(n2236), .Y(n2235) );
  OAI22XL U13890 ( .A0(n8175), .A1(n9324), .B0(n8171), .B1(n9322), .Y(n2236)
         );
  AOI221XL U13891 ( .A0(\xArray[13][10] ), .A1(n8180), .B0(\xArray[1][10] ), 
        .B1(n8178), .C0(n2227), .Y(n2226) );
  OAI22XL U13892 ( .A0(n8175), .A1(n9316), .B0(n8171), .B1(n9314), .Y(n2227)
         );
  AOI221XL U13893 ( .A0(\xArray[13][11] ), .A1(n8180), .B0(\xArray[1][11] ), 
        .B1(n8178), .C0(n2218), .Y(n2217) );
  OA22X1 U13894 ( .A0(n8322), .A1(n1506), .B0(n7728), .B1(n1709), .Y(n2216) );
  OAI22XL U13895 ( .A0(n8175), .A1(n9308), .B0(n8171), .B1(n9306), .Y(n2218)
         );
  OAI221X1 U13896 ( .A0(\xArray[7][17] ), .A1(n8296), .B0(\xArray[11][17] ), 
        .B1(n8242), .C0(n1209), .Y(n637) );
  AOI2BB2X1 U13897 ( .B0(n9256), .B1(n8212), .A0N(\xArray[15][17] ), .A1N(
        n8255), .Y(n1209) );
  OAI221X1 U13898 ( .A0(\xArray[7][18] ), .A1(n8297), .B0(\xArray[11][18] ), 
        .B1(n8243), .C0(n1204), .Y(n629) );
  OAI221X1 U13899 ( .A0(\xArray[4][18] ), .A1(n8286), .B0(\xArray[8][18] ), 
        .B1(n8232), .C0(n2161), .Y(n1476) );
  OA22X1 U13900 ( .A0(\xArray[0][18] ), .A1(n8191), .B0(\xArray[12][18] ), 
        .B1(n8265), .Y(n2161) );
  OAI221X1 U13901 ( .A0(\xArray[4][19] ), .A1(n8286), .B0(\xArray[8][19] ), 
        .B1(n8232), .C0(n2152), .Y(n1472) );
  OA22X1 U13902 ( .A0(\xArray[0][19] ), .A1(n8191), .B0(\xArray[12][19] ), 
        .B1(n8265), .Y(n2152) );
  OAI221X1 U13903 ( .A0(\xArray[8][17] ), .A1(n8297), .B0(\xArray[12][17] ), 
        .B1(n8243), .C0(n1208), .Y(n639) );
  OA22X1 U13904 ( .A0(\xArray[4][17] ), .A1(n8198), .B0(\xArray[0][17] ), .B1(
        n8267), .Y(n1208) );
  OAI221X1 U13905 ( .A0(\xArray[8][18] ), .A1(n8297), .B0(\xArray[12][18] ), 
        .B1(n8243), .C0(n1203), .Y(n631) );
  OAI221X1 U13906 ( .A0(\xArray[6][18] ), .A1(n8293), .B0(\xArray[10][18] ), 
        .B1(n8239), .C0(n1479), .Y(n920) );
  OAI221X1 U13907 ( .A0(\xArray[3][18] ), .A1(n8286), .B0(\xArray[7][18] ), 
        .B1(n8232), .C0(n2160), .Y(n1478) );
  OA22X1 U13908 ( .A0(\xArray[15][18] ), .A1(n8191), .B0(\xArray[11][18] ), 
        .B1(n8265), .Y(n2160) );
  OAI221X1 U13909 ( .A0(\xArray[3][19] ), .A1(n8286), .B0(\xArray[7][19] ), 
        .B1(n8232), .C0(n2151), .Y(n1474) );
  OA22X1 U13910 ( .A0(\xArray[15][19] ), .A1(n8191), .B0(\xArray[11][19] ), 
        .B1(n8265), .Y(n2151) );
  OAI221X1 U13911 ( .A0(\xArray[5][18] ), .A1(n8281), .B0(\xArray[9][18] ), 
        .B1(n8227), .C0(n1689), .Y(n1202) );
  OA22X1 U13912 ( .A0(\xArray[1][18] ), .A1(n8188), .B0(\xArray[13][18] ), 
        .B1(n8259), .Y(n1689) );
  OAI221X1 U13913 ( .A0(\xArray[5][19] ), .A1(n8281), .B0(\xArray[9][19] ), 
        .B1(n8227), .C0(n1686), .Y(n1197) );
  OAI221XL U13914 ( .A0(\xArray[9][17] ), .A1(n8290), .B0(\xArray[13][17] ), 
        .B1(n8236), .C0(n924), .Y(n638) );
  OA22X1 U13915 ( .A0(\xArray[5][17] ), .A1(n8195), .B0(\xArray[1][17] ), .B1(
        n8269), .Y(n924) );
  OAI221XL U13916 ( .A0(\xArray[9][18] ), .A1(n8290), .B0(\xArray[13][18] ), 
        .B1(n8236), .C0(n921), .Y(n630) );
  OA22X1 U13917 ( .A0(\xArray[5][18] ), .A1(n8195), .B0(\xArray[1][18] ), .B1(
        n8269), .Y(n921) );
  OAI221XL U13918 ( .A0(\xArray[2][15] ), .A1(n8285), .B0(\xArray[6][15] ), 
        .B1(n8231), .C0(n2185), .Y(n1697) );
  OAI221XL U13919 ( .A0(\xArray[2][16] ), .A1(n8285), .B0(\xArray[6][16] ), 
        .B1(n8231), .C0(n2176), .Y(n1694) );
  OAI222XL U13920 ( .A0(n717), .A1(n8340), .B0(n718), .B1(n8308), .C0(n719), 
        .C1(n7712), .Y(n712) );
  AOI221XL U13921 ( .A0(\xArray[14][7] ), .A1(n6573), .B0(\xArray[2][7] ), 
        .B1(n8361), .C0(n714), .Y(n713) );
  OAI22XL U13922 ( .A0(n8357), .A1(n9339), .B0(n8355), .B1(n9341), .Y(n714) );
  OAI222XL U13923 ( .A0(n725), .A1(n8340), .B0(n726), .B1(n8308), .C0(n727), 
        .C1(n7712), .Y(n720) );
  AOI221XL U13924 ( .A0(\xArray[14][6] ), .A1(n6573), .B0(\xArray[2][6] ), 
        .B1(n8361), .C0(n722), .Y(n721) );
  OAI22XL U13925 ( .A0(n8357), .A1(n9347), .B0(n8355), .B1(n9349), .Y(n722) );
  OAI222XL U13926 ( .A0(n733), .A1(n8340), .B0(n734), .B1(n8308), .C0(n735), 
        .C1(n7712), .Y(n728) );
  AOI221XL U13927 ( .A0(\xArray[14][5] ), .A1(n6573), .B0(\xArray[2][5] ), 
        .B1(n8361), .C0(n730), .Y(n729) );
  OAI22XL U13928 ( .A0(n8359), .A1(n9355), .B0(n8355), .B1(n9357), .Y(n730) );
  OAI222XL U13929 ( .A0(n741), .A1(n8340), .B0(n742), .B1(n8308), .C0(n743), 
        .C1(n7712), .Y(n736) );
  AOI221XL U13930 ( .A0(\xArray[14][4] ), .A1(n6573), .B0(\xArray[2][4] ), 
        .B1(n8361), .C0(n738), .Y(n737) );
  OAI22XL U13931 ( .A0(n8359), .A1(n9363), .B0(n8355), .B1(n9365), .Y(n738) );
  OAI221XL U13932 ( .A0(n7424), .A1(n8065), .B0(n7539), .B1(n8062), .C0(n3193), 
        .Y(N28281) );
  OAI221XL U13933 ( .A0(n7424), .A1(n8142), .B0(n7539), .B1(n8139), .C0(n2678), 
        .Y(N28665) );
  OAI221XL U13934 ( .A0(n7426), .A1(n8065), .B0(n7538), .B1(n8061), .C0(n3192), 
        .Y(N28282) );
  OAI221XL U13935 ( .A0(n7426), .A1(n8142), .B0(n7538), .B1(n8140), .C0(n2676), 
        .Y(N28666) );
  OAI221XL U13936 ( .A0(n7428), .A1(n8066), .B0(n7537), .B1(n8063), .C0(n3191), 
        .Y(N28283) );
  OAI221XL U13937 ( .A0(n7428), .A1(n8143), .B0(n7537), .B1(n8140), .C0(n2674), 
        .Y(N28667) );
  OAI221XL U13938 ( .A0(n7430), .A1(n8066), .B0(n7536), .B1(n8063), .C0(n3190), 
        .Y(N28284) );
  OAI221XL U13939 ( .A0(n7430), .A1(n8143), .B0(n7536), .B1(n8138), .C0(n2672), 
        .Y(N28668) );
  OAI221XL U13940 ( .A0(n7432), .A1(n8066), .B0(n7535), .B1(n8063), .C0(n3189), 
        .Y(N28285) );
  OAI221XL U13941 ( .A0(n7432), .A1(n8143), .B0(n7535), .B1(n8138), .C0(n2670), 
        .Y(N28669) );
  AND4X1 U13942 ( .A(n4389), .B(n4390), .C(n4391), .D(n4392), .Y(n2448) );
  AOI221XL U13943 ( .A0(n7963), .A1(\xArray[9][24] ), .B0(\xArray[8][24] ), 
        .B1(n7961), .C0(n4393), .Y(n4392) );
  AOI221XL U13944 ( .A0(n7949), .A1(n7423), .B0(n7946), .B1(\xArray[2][24] ), 
        .C0(n4395), .Y(n4391) );
  AND4X1 U13945 ( .A(n4371), .B(n4372), .C(n4373), .D(n4374), .Y(n2445) );
  AOI221XL U13946 ( .A0(n7964), .A1(\xArray[9][25] ), .B0(\xArray[8][25] ), 
        .B1(n7961), .C0(n4375), .Y(n4374) );
  AOI221XL U13947 ( .A0(n7949), .A1(n7425), .B0(n7946), .B1(\xArray[2][25] ), 
        .C0(n4377), .Y(n4373) );
  AND4X1 U13948 ( .A(n4353), .B(n4354), .C(n4355), .D(n4356), .Y(n2442) );
  AOI221XL U13949 ( .A0(n7963), .A1(\xArray[9][26] ), .B0(\xArray[8][26] ), 
        .B1(n7961), .C0(n4357), .Y(n4356) );
  AOI221XL U13950 ( .A0(n7949), .A1(n7427), .B0(n7946), .B1(\xArray[2][26] ), 
        .C0(n4359), .Y(n4355) );
  AND4X1 U13951 ( .A(n4335), .B(n4336), .C(n4337), .D(n4338), .Y(n2439) );
  AOI221XL U13952 ( .A0(n7964), .A1(\xArray[9][27] ), .B0(\xArray[8][27] ), 
        .B1(n7960), .C0(n4339), .Y(n4338) );
  AOI221XL U13953 ( .A0(n7949), .A1(n7429), .B0(n7946), .B1(\xArray[2][27] ), 
        .C0(n4341), .Y(n4337) );
  OAI221X1 U13954 ( .A0(\xArray[7][19] ), .A1(n8297), .B0(\xArray[11][19] ), 
        .B1(n8243), .C0(n1199), .Y(n621) );
  OAI221X1 U13955 ( .A0(\xArray[7][20] ), .A1(n8297), .B0(\xArray[11][20] ), 
        .B1(n8243), .C0(n1194), .Y(n613) );
  OAI221X1 U13956 ( .A0(\xArray[4][20] ), .A1(n8286), .B0(\xArray[8][20] ), 
        .B1(n8232), .C0(n2143), .Y(n1468) );
  OA22X1 U13957 ( .A0(\xArray[0][20] ), .A1(n8191), .B0(\xArray[12][20] ), 
        .B1(n8265), .Y(n2143) );
  OAI221X1 U13958 ( .A0(\xArray[4][21] ), .A1(n8286), .B0(\xArray[8][21] ), 
        .B1(n8232), .C0(n2134), .Y(n1464) );
  OA22X1 U13959 ( .A0(\xArray[0][21] ), .A1(n8191), .B0(\xArray[12][21] ), 
        .B1(n8266), .Y(n2134) );
  OAI221X1 U13960 ( .A0(\xArray[8][19] ), .A1(n8297), .B0(\xArray[12][19] ), 
        .B1(n8243), .C0(n1198), .Y(n623) );
  OAI221X1 U13961 ( .A0(\xArray[8][20] ), .A1(n8297), .B0(\xArray[12][20] ), 
        .B1(n8243), .C0(n1193), .Y(n615) );
  OAI221X1 U13962 ( .A0(\xArray[6][19] ), .A1(n8293), .B0(\xArray[10][19] ), 
        .B1(n8239), .C0(n1475), .Y(n917) );
  OAI221X1 U13963 ( .A0(\xArray[6][20] ), .A1(n8293), .B0(\xArray[10][20] ), 
        .B1(n8239), .C0(n1471), .Y(n914) );
  OAI221X1 U13964 ( .A0(\xArray[3][20] ), .A1(n8286), .B0(\xArray[7][20] ), 
        .B1(n8232), .C0(n2142), .Y(n1470) );
  OA22X1 U13965 ( .A0(\xArray[15][20] ), .A1(n8191), .B0(\xArray[11][20] ), 
        .B1(n8265), .Y(n2142) );
  OAI221X1 U13966 ( .A0(\xArray[5][20] ), .A1(n8281), .B0(\xArray[9][20] ), 
        .B1(n8227), .C0(n1683), .Y(n1192) );
  OAI221X1 U13967 ( .A0(\xArray[5][21] ), .A1(n8281), .B0(\xArray[9][21] ), 
        .B1(n8227), .C0(n1680), .Y(n1187) );
  OAI221XL U13968 ( .A0(\xArray[9][19] ), .A1(n8291), .B0(\xArray[13][19] ), 
        .B1(n8237), .C0(n918), .Y(n622) );
  OA22X1 U13969 ( .A0(\xArray[5][19] ), .A1(n8195), .B0(\xArray[1][19] ), .B1(
        n8269), .Y(n918) );
  OAI221XL U13970 ( .A0(\xArray[9][20] ), .A1(n8291), .B0(\xArray[13][20] ), 
        .B1(n8237), .C0(n915), .Y(n614) );
  OAI221XL U13971 ( .A0(\xArray[2][17] ), .A1(n8286), .B0(\xArray[6][17] ), 
        .B1(n8232), .C0(n2167), .Y(n1691) );
  OAI221XL U13972 ( .A0(\xArray[2][18] ), .A1(n8286), .B0(\xArray[6][18] ), 
        .B1(n8232), .C0(n2158), .Y(n1688) );
  AOI221XL U13973 ( .A0(n7949), .A1(n7417), .B0(n7946), .B1(\xArray[2][21] ), 
        .C0(n4449), .Y(n4445) );
  OAI222XL U13974 ( .A0(n9226), .A1(n7942), .B0(n8658), .B1(n7940), .C0(n7937), 
        .C1(n9225), .Y(n4449) );
  AOI221XL U13975 ( .A0(n7949), .A1(n7419), .B0(n7946), .B1(\xArray[2][22] ), 
        .C0(n4431), .Y(n4427) );
  OAI222XL U13976 ( .A0(n9218), .A1(n7942), .B0(n8653), .B1(n7940), .C0(n7937), 
        .C1(n9217), .Y(n4431) );
  OAI221XL U13977 ( .A0(n7418), .A1(n8065), .B0(n7542), .B1(n8062), .C0(n3196), 
        .Y(N28278) );
  OAI221XL U13978 ( .A0(n7418), .A1(n8142), .B0(n7542), .B1(n8138), .C0(n2684), 
        .Y(N28662) );
  OAI221XL U13979 ( .A0(n7420), .A1(n8065), .B0(n7541), .B1(n8062), .C0(n3195), 
        .Y(N28279) );
  OAI221XL U13980 ( .A0(n7420), .A1(n8142), .B0(n7541), .B1(n8139), .C0(n2682), 
        .Y(N28663) );
  OAI221XL U13981 ( .A0(n7422), .A1(n8065), .B0(n7540), .B1(n8062), .C0(n3194), 
        .Y(N28280) );
  OAI221XL U13982 ( .A0(n7422), .A1(n8142), .B0(n7540), .B1(n8139), .C0(n2680), 
        .Y(N28664) );
  AND4X1 U13983 ( .A(n4443), .B(n4444), .C(n4445), .D(n4446), .Y(n2457) );
  AOI221XL U13984 ( .A0(n7963), .A1(\xArray[9][21] ), .B0(\xArray[8][21] ), 
        .B1(n7961), .C0(n4447), .Y(n4446) );
  AOI221XL U13985 ( .A0(n8661), .A1(n7993), .B0(n8662), .B1(n8030), .C0(n4452), 
        .Y(n4444) );
  AND4X1 U13986 ( .A(n4425), .B(n4426), .C(n4427), .D(n4428), .Y(n2454) );
  AOI221XL U13987 ( .A0(n7964), .A1(\xArray[9][22] ), .B0(\xArray[8][22] ), 
        .B1(n7961), .C0(n4429), .Y(n4428) );
  AOI221XL U13988 ( .A0(n8656), .A1(n7993), .B0(n8657), .B1(n8030), .C0(n4434), 
        .Y(n4426) );
  AND4X1 U13989 ( .A(n4407), .B(n4408), .C(n4409), .D(n4410), .Y(n2451) );
  AOI221XL U13990 ( .A0(n7964), .A1(\xArray[9][23] ), .B0(\xArray[8][23] ), 
        .B1(n7960), .C0(n4411), .Y(n4410) );
  AOI221XL U13991 ( .A0(n7949), .A1(n7421), .B0(n7946), .B1(\xArray[2][23] ), 
        .C0(n4413), .Y(n4409) );
  MX4X1 U13992 ( .A(\bArray[12][16] ), .B(\bArray[13][16] ), .C(
        \bArray[14][16] ), .D(\bArray[15][16] ), .S0(n7205), .S1(n7217), .Y(
        n7008) );
  MX4X1 U13993 ( .A(\bArray[8][16] ), .B(\bArray[9][16] ), .C(\bArray[10][16] ), .D(\bArray[11][16] ), .S0(n7205), .S1(n7217), .Y(n7009) );
  MX4X1 U13994 ( .A(\bArray[4][16] ), .B(\bArray[5][16] ), .C(\bArray[6][16] ), 
        .D(\bArray[7][16] ), .S0(n7205), .S1(n7217), .Y(n7010) );
  AOI221XL U13995 ( .A0(\xArray[13][12] ), .A1(n8180), .B0(\xArray[1][12] ), 
        .B1(n8178), .C0(n2209), .Y(n2208) );
  OA22X1 U13996 ( .A0(n8322), .A1(n1502), .B0(n7728), .B1(n1706), .Y(n2207) );
  OAI22XL U13997 ( .A0(n8175), .A1(n9300), .B0(n8172), .B1(n9298), .Y(n2209)
         );
  AOI221XL U13998 ( .A0(\xArray[13][13] ), .A1(n8180), .B0(\xArray[1][13] ), 
        .B1(n8178), .C0(n2200), .Y(n2199) );
  OA22X1 U13999 ( .A0(n8322), .A1(n1498), .B0(n7730), .B1(n1703), .Y(n2198) );
  OAI22XL U14000 ( .A0(n8173), .A1(n9292), .B0(n8172), .B1(n9290), .Y(n2200)
         );
  AOI221XL U14001 ( .A0(\xArray[13][14] ), .A1(n8180), .B0(\xArray[1][14] ), 
        .B1(n8178), .C0(n2191), .Y(n2190) );
  OA22X1 U14002 ( .A0(n8322), .A1(n1494), .B0(n7728), .B1(n1700), .Y(n2189) );
  OAI22XL U14003 ( .A0(n8175), .A1(n9284), .B0(n8172), .B1(n9282), .Y(n2191)
         );
  AOI221XL U14004 ( .A0(\xArray[13][15] ), .A1(n8180), .B0(\xArray[1][15] ), 
        .B1(n8178), .C0(n2182), .Y(n2181) );
  OA22X1 U14005 ( .A0(n8322), .A1(n1490), .B0(n7728), .B1(n1697), .Y(n2180) );
  OAI22XL U14006 ( .A0(n8173), .A1(n9276), .B0(n8172), .B1(n9274), .Y(n2182)
         );
  OAI221X1 U14007 ( .A0(\xArray[7][21] ), .A1(n8297), .B0(\xArray[11][21] ), 
        .B1(n8243), .C0(n1189), .Y(n605) );
  OAI221X1 U14008 ( .A0(\xArray[7][22] ), .A1(n8297), .B0(\xArray[11][22] ), 
        .B1(n8243), .C0(n1184), .Y(n597) );
  OAI221X1 U14009 ( .A0(\xArray[4][22] ), .A1(n8286), .B0(\xArray[8][22] ), 
        .B1(n8232), .C0(n2125), .Y(n1460) );
  OA22X1 U14010 ( .A0(\xArray[0][22] ), .A1(n8191), .B0(\xArray[12][22] ), 
        .B1(n8266), .Y(n2125) );
  OAI221X1 U14011 ( .A0(\xArray[4][23] ), .A1(n8287), .B0(\xArray[8][23] ), 
        .B1(n8233), .C0(n2116), .Y(n1456) );
  OA22X1 U14012 ( .A0(\xArray[0][23] ), .A1(n8191), .B0(\xArray[12][23] ), 
        .B1(n8266), .Y(n2116) );
  OAI221X1 U14013 ( .A0(\xArray[8][21] ), .A1(n8297), .B0(\xArray[12][21] ), 
        .B1(n8243), .C0(n1188), .Y(n607) );
  OAI221X1 U14014 ( .A0(\xArray[8][22] ), .A1(n8297), .B0(\xArray[12][22] ), 
        .B1(n8243), .C0(n1183), .Y(n599) );
  OAI221X1 U14015 ( .A0(\xArray[6][21] ), .A1(n8293), .B0(\xArray[10][21] ), 
        .B1(n8239), .C0(n1467), .Y(n911) );
  OAI221X1 U14016 ( .A0(\xArray[3][21] ), .A1(n8286), .B0(\xArray[7][21] ), 
        .B1(n8232), .C0(n2133), .Y(n1466) );
  OA22X1 U14017 ( .A0(\xArray[15][21] ), .A1(n8191), .B0(\xArray[11][21] ), 
        .B1(n8266), .Y(n2133) );
  OAI221X1 U14018 ( .A0(\xArray[6][22] ), .A1(n8293), .B0(\xArray[10][22] ), 
        .B1(n8239), .C0(n1463), .Y(n908) );
  OAI221X1 U14019 ( .A0(\xArray[3][22] ), .A1(n8286), .B0(\xArray[7][22] ), 
        .B1(n8232), .C0(n2124), .Y(n1462) );
  OA22X1 U14020 ( .A0(\xArray[15][22] ), .A1(n8191), .B0(\xArray[11][22] ), 
        .B1(n8266), .Y(n2124) );
  OAI221X1 U14021 ( .A0(\xArray[5][22] ), .A1(n8281), .B0(\xArray[9][22] ), 
        .B1(n8227), .C0(n1677), .Y(n1182) );
  OAI221X1 U14022 ( .A0(\xArray[5][23] ), .A1(n8282), .B0(\xArray[9][23] ), 
        .B1(n8228), .C0(n1674), .Y(n1177) );
  OA22X1 U14023 ( .A0(\xArray[1][23] ), .A1(n8188), .B0(\xArray[13][23] ), 
        .B1(n8261), .Y(n1674) );
  OAI221XL U14024 ( .A0(\xArray[9][21] ), .A1(n8291), .B0(\xArray[13][21] ), 
        .B1(n8237), .C0(n912), .Y(n606) );
  OAI221XL U14025 ( .A0(\xArray[2][19] ), .A1(n8286), .B0(\xArray[6][19] ), 
        .B1(n8232), .C0(n2149), .Y(n1685) );
  OAI221XL U14026 ( .A0(\xArray[2][20] ), .A1(n8286), .B0(\xArray[6][20] ), 
        .B1(n8232), .C0(n2140), .Y(n1682) );
  OAI222XL U14027 ( .A0(n685), .A1(n8340), .B0(n686), .B1(n8308), .C0(n687), 
        .C1(n7712), .Y(n680) );
  AOI221XL U14028 ( .A0(\xArray[14][11] ), .A1(n6573), .B0(\xArray[2][11] ), 
        .B1(n8361), .C0(n682), .Y(n681) );
  OAI22XL U14029 ( .A0(n8357), .A1(n9307), .B0(n8355), .B1(n9309), .Y(n682) );
  OAI222XL U14030 ( .A0(n693), .A1(n8340), .B0(n694), .B1(n8308), .C0(n695), 
        .C1(n7712), .Y(n688) );
  AOI221XL U14031 ( .A0(\xArray[14][10] ), .A1(n6573), .B0(\xArray[2][10] ), 
        .B1(n8361), .C0(n690), .Y(n689) );
  OAI22XL U14032 ( .A0(n8357), .A1(n9315), .B0(n8355), .B1(n9317), .Y(n690) );
  OAI222XL U14033 ( .A0(n701), .A1(n8340), .B0(n702), .B1(n8308), .C0(n703), 
        .C1(n7712), .Y(n696) );
  AOI221XL U14034 ( .A0(\xArray[14][9] ), .A1(n6573), .B0(\xArray[2][9] ), 
        .B1(n8361), .C0(n698), .Y(n697) );
  OAI22XL U14035 ( .A0(n8357), .A1(n9323), .B0(n8355), .B1(n9325), .Y(n698) );
  OAI222XL U14036 ( .A0(n709), .A1(n8340), .B0(n710), .B1(n8308), .C0(n711), 
        .C1(n7712), .Y(n704) );
  AOI221XL U14037 ( .A0(\xArray[14][8] ), .A1(n6573), .B0(\xArray[2][8] ), 
        .B1(n8361), .C0(n706), .Y(n705) );
  OAI22XL U14038 ( .A0(n8357), .A1(n9331), .B0(n8355), .B1(n9333), .Y(n706) );
  OAI221XL U14039 ( .A0(n7408), .A1(n8065), .B0(n7547), .B1(n8061), .C0(n3201), 
        .Y(N28273) );
  OAI221XL U14040 ( .A0(n7408), .A1(n8142), .B0(n7547), .B1(n8138), .C0(n2694), 
        .Y(N28657) );
  OAI221XL U14041 ( .A0(n7410), .A1(n8065), .B0(n7546), .B1(n8061), .C0(n3200), 
        .Y(N28274) );
  OAI221XL U14042 ( .A0(n7410), .A1(n8142), .B0(n7546), .B1(n8138), .C0(n2692), 
        .Y(N28658) );
  OAI221XL U14043 ( .A0(n7412), .A1(n8065), .B0(n7545), .B1(n8061), .C0(n3199), 
        .Y(N28275) );
  OAI221XL U14044 ( .A0(n7412), .A1(n8142), .B0(n7545), .B1(n8138), .C0(n2690), 
        .Y(N28659) );
  OAI221XL U14045 ( .A0(n7414), .A1(n8065), .B0(n7544), .B1(n8061), .C0(n3198), 
        .Y(N28276) );
  OAI221XL U14046 ( .A0(n7414), .A1(n8142), .B0(n7544), .B1(n8138), .C0(n2688), 
        .Y(N28660) );
  OAI221XL U14047 ( .A0(n7416), .A1(n8065), .B0(n7543), .B1(n8061), .C0(n3197), 
        .Y(N28277) );
  OAI221XL U14048 ( .A0(n7416), .A1(n8142), .B0(n7543), .B1(n8138), .C0(n2686), 
        .Y(N28661) );
  MX4X1 U14049 ( .A(n6792), .B(n6790), .C(n6791), .D(n6789), .S0(n7005), .S1(
        n7003), .Y(N25583) );
  MX4X1 U14050 ( .A(n6788), .B(n6786), .C(n6787), .D(n6785), .S0(n7005), .S1(
        n7003), .Y(N25584) );
  MX4X1 U14051 ( .A(\bArray[0][16] ), .B(\bArray[1][16] ), .C(\bArray[2][16] ), 
        .D(\bArray[3][16] ), .S0(n7205), .S1(n7217), .Y(n7011) );
  CLKBUFX3 U14052 ( .A(n2475), .Y(n7406) );
  AND4X1 U14053 ( .A(n4551), .B(n4552), .C(n4553), .D(n4554), .Y(n2475) );
  AOI221XL U14054 ( .A0(n7964), .A1(\xArray[9][15] ), .B0(\xArray[8][15] ), 
        .B1(n7959), .C0(n4555), .Y(n4554) );
  AOI221XL U14055 ( .A0(n6603), .A1(n7405), .B0(n7944), .B1(\xArray[2][15] ), 
        .C0(n4557), .Y(n4553) );
  AND4X1 U14056 ( .A(n4533), .B(n4534), .C(n4535), .D(n4536), .Y(n2472) );
  AOI221XL U14057 ( .A0(n7965), .A1(\xArray[9][16] ), .B0(\xArray[8][16] ), 
        .B1(n7960), .C0(n4537), .Y(n4536) );
  AOI221XL U14058 ( .A0(n7949), .A1(n7407), .B0(n7946), .B1(\xArray[2][16] ), 
        .C0(n4539), .Y(n4535) );
  AND4X1 U14059 ( .A(n4515), .B(n4516), .C(n4517), .D(n4518), .Y(n2469) );
  AOI221XL U14060 ( .A0(n7962), .A1(\xArray[9][17] ), .B0(\xArray[8][17] ), 
        .B1(n7959), .C0(n4519), .Y(n4518) );
  AOI221XL U14061 ( .A0(n7949), .A1(n7409), .B0(n7946), .B1(\xArray[2][17] ), 
        .C0(n4521), .Y(n4517) );
  AND4X1 U14062 ( .A(n4497), .B(n4498), .C(n4499), .D(n4500), .Y(n2466) );
  AOI221XL U14063 ( .A0(n7964), .A1(\xArray[9][18] ), .B0(\xArray[8][18] ), 
        .B1(n7961), .C0(n4501), .Y(n4500) );
  AOI221XL U14064 ( .A0(n7949), .A1(n7411), .B0(n7946), .B1(\xArray[2][18] ), 
        .C0(n4503), .Y(n4499) );
  AND4X1 U14065 ( .A(n4479), .B(n4480), .C(n4481), .D(n4482), .Y(n2463) );
  AOI221XL U14066 ( .A0(n3659), .A1(\xArray[9][19] ), .B0(\xArray[8][19] ), 
        .B1(n7960), .C0(n4483), .Y(n4482) );
  AOI221XL U14067 ( .A0(n7949), .A1(n7413), .B0(n7946), .B1(\xArray[2][19] ), 
        .C0(n4485), .Y(n4481) );
  AND4X1 U14068 ( .A(n4461), .B(n4462), .C(n4463), .D(n4464), .Y(n2460) );
  AOI221XL U14069 ( .A0(n7963), .A1(\xArray[9][20] ), .B0(\xArray[8][20] ), 
        .B1(n7961), .C0(n4465), .Y(n4464) );
  AOI221XL U14070 ( .A0(n7949), .A1(n7415), .B0(n7946), .B1(\xArray[2][20] ), 
        .C0(n4467), .Y(n4463) );
  CLKBUFX3 U14071 ( .A(N1762), .Y(n8409) );
  CLKBUFX3 U14072 ( .A(N1761), .Y(n8410) );
  CLKBUFX3 U14073 ( .A(N1757), .Y(n8414) );
  MX4X1 U14074 ( .A(\bArray[4][18] ), .B(\bArray[5][18] ), .C(\bArray[6][18] ), 
        .D(\bArray[7][18] ), .S0(n7206), .S1(n7218), .Y(n7018) );
  OAI221X1 U14075 ( .A0(\xArray[7][24] ), .A1(n8297), .B0(\xArray[11][24] ), 
        .B1(n8243), .C0(n1174), .Y(n581) );
  OAI221X1 U14076 ( .A0(\xArray[4][24] ), .A1(n8287), .B0(\xArray[8][24] ), 
        .B1(n8233), .C0(n2107), .Y(n1452) );
  OAI221X1 U14077 ( .A0(\xArray[4][25] ), .A1(n8287), .B0(\xArray[8][25] ), 
        .B1(n8233), .C0(n2098), .Y(n1448) );
  OAI221X1 U14078 ( .A0(\xArray[8][23] ), .A1(n8297), .B0(\xArray[12][23] ), 
        .B1(n8243), .C0(n1178), .Y(n591) );
  OAI221X1 U14079 ( .A0(\xArray[8][24] ), .A1(n8297), .B0(\xArray[12][24] ), 
        .B1(n8243), .C0(n1173), .Y(n583) );
  OAI221X1 U14080 ( .A0(\xArray[6][23] ), .A1(n8293), .B0(\xArray[10][23] ), 
        .B1(n8239), .C0(n1459), .Y(n905) );
  OAI221X1 U14081 ( .A0(\xArray[3][23] ), .A1(n8287), .B0(\xArray[7][23] ), 
        .B1(n8233), .C0(n2115), .Y(n1458) );
  OA22X1 U14082 ( .A0(\xArray[15][23] ), .A1(n8191), .B0(\xArray[11][23] ), 
        .B1(n8266), .Y(n2115) );
  OAI221X1 U14083 ( .A0(\xArray[6][24] ), .A1(n8293), .B0(\xArray[10][24] ), 
        .B1(n8239), .C0(n1455), .Y(n902) );
  OAI221X1 U14084 ( .A0(\xArray[3][24] ), .A1(n8287), .B0(\xArray[7][24] ), 
        .B1(n8233), .C0(n2106), .Y(n1454) );
  OAI221X1 U14085 ( .A0(\xArray[5][24] ), .A1(n8282), .B0(\xArray[9][24] ), 
        .B1(n8228), .C0(n1671), .Y(n1172) );
  OAI221X1 U14086 ( .A0(\xArray[5][25] ), .A1(n8282), .B0(\xArray[9][25] ), 
        .B1(n8228), .C0(n1668), .Y(n1167) );
  OAI221XL U14087 ( .A0(\xArray[9][22] ), .A1(n8291), .B0(\xArray[13][22] ), 
        .B1(n8237), .C0(n909), .Y(n598) );
  OAI221XL U14088 ( .A0(\xArray[9][23] ), .A1(n8291), .B0(\xArray[13][23] ), 
        .B1(n8237), .C0(n906), .Y(n590) );
  OAI221XL U14089 ( .A0(\xArray[2][22] ), .A1(n8287), .B0(\xArray[6][22] ), 
        .B1(n8233), .C0(n2122), .Y(n1676) );
  OAI222XL U14090 ( .A0(n677), .A1(n8339), .B0(n678), .B1(n8307), .C0(n679), 
        .C1(n7713), .Y(n672) );
  AOI221XL U14091 ( .A0(\xArray[14][12] ), .A1(n6573), .B0(\xArray[2][12] ), 
        .B1(n8361), .C0(n674), .Y(n673) );
  OAI22XL U14092 ( .A0(n8359), .A1(n9299), .B0(n8353), .B1(n9301), .Y(n674) );
  AOI221XL U14093 ( .A0(n7947), .A1(n7399), .B0(n7946), .B1(\xArray[2][12] ), 
        .C0(n4611), .Y(n4607) );
  OAI222XL U14094 ( .A0(n9298), .A1(n7943), .B0(n8703), .B1(n7939), .C0(n3671), 
        .C1(n9297), .Y(n4611) );
  OAI221XL U14095 ( .A0(n7400), .A1(n8065), .B0(n7551), .B1(n8061), .C0(n3205), 
        .Y(N28269) );
  OAI221XL U14096 ( .A0(n7400), .A1(n8142), .B0(n7551), .B1(n8138), .C0(n2702), 
        .Y(N28653) );
  OAI221XL U14097 ( .A0(n7402), .A1(n8065), .B0(n7550), .B1(n8061), .C0(n3204), 
        .Y(N28270) );
  OAI221XL U14098 ( .A0(n7402), .A1(n8142), .B0(n7550), .B1(n8138), .C0(n2700), 
        .Y(N28654) );
  OAI221XL U14099 ( .A0(n7404), .A1(n8065), .B0(n7549), .B1(n8061), .C0(n3203), 
        .Y(N28271) );
  OAI221XL U14100 ( .A0(n7404), .A1(n8142), .B0(n7549), .B1(n8138), .C0(n2698), 
        .Y(N28655) );
  OAI221XL U14101 ( .A0(n7406), .A1(n8065), .B0(n7548), .B1(n8061), .C0(n3202), 
        .Y(N28272) );
  OAI221XL U14102 ( .A0(n7406), .A1(n8142), .B0(n7548), .B1(n8138), .C0(n2696), 
        .Y(N28656) );
  MX4X1 U14103 ( .A(n6800), .B(n6798), .C(n6799), .D(n6797), .S0(n7005), .S1(
        n7003), .Y(N25581) );
  MX4X1 U14104 ( .A(n6796), .B(n6794), .C(n6795), .D(n6793), .S0(n7005), .S1(
        n7003), .Y(N25582) );
  OAI221XL U14105 ( .A0(\xArray[2][21] ), .A1(n8286), .B0(\xArray[6][21] ), 
        .B1(n8232), .C0(n2131), .Y(n1679) );
  MX4X1 U14106 ( .A(\bArray[0][18] ), .B(\bArray[1][18] ), .C(\bArray[2][18] ), 
        .D(\bArray[3][18] ), .S0(n7206), .S1(n7218), .Y(n7019) );
  AND4X1 U14107 ( .A(n4605), .B(n4606), .C(n4607), .D(n4608), .Y(n2484) );
  AOI221XL U14108 ( .A0(n7965), .A1(\xArray[9][12] ), .B0(\xArray[8][12] ), 
        .B1(n7959), .C0(n4609), .Y(n4608) );
  AOI221XL U14109 ( .A0(n8706), .A1(n7992), .B0(n8707), .B1(n8029), .C0(n4614), 
        .Y(n4606) );
  AND4X1 U14110 ( .A(n4587), .B(n4588), .C(n4589), .D(n4590), .Y(n2481) );
  AOI221XL U14111 ( .A0(n7962), .A1(\xArray[9][13] ), .B0(\xArray[8][13] ), 
        .B1(n7960), .C0(n4591), .Y(n4590) );
  AOI221XL U14112 ( .A0(n7949), .A1(n7401), .B0(n7944), .B1(\xArray[2][13] ), 
        .C0(n4593), .Y(n4589) );
  AND4X1 U14113 ( .A(n4569), .B(n4570), .C(n4571), .D(n4572), .Y(n2478) );
  AOI221XL U14114 ( .A0(n7964), .A1(\xArray[9][14] ), .B0(\xArray[8][14] ), 
        .B1(n7960), .C0(n4573), .Y(n4572) );
  AOI221XL U14115 ( .A0(n7948), .A1(n7403), .B0(n7944), .B1(\xArray[2][14] ), 
        .C0(n4575), .Y(n4571) );
  CLKBUFX3 U14116 ( .A(N1764), .Y(n8407) );
  CLKBUFX3 U14117 ( .A(N1763), .Y(n8408) );
  CLKBUFX3 U14118 ( .A(N1760), .Y(n8411) );
  CLKBUFX3 U14119 ( .A(N1759), .Y(n8412) );
  CLKBUFX3 U14120 ( .A(N1758), .Y(n8413) );
  AOI221XL U14121 ( .A0(\xArray[13][16] ), .A1(n8181), .B0(\xArray[1][16] ), 
        .B1(n8177), .C0(n2173), .Y(n2172) );
  OAI22XL U14122 ( .A0(n8173), .A1(n9268), .B0(n8172), .B1(n9266), .Y(n2173)
         );
  AOI221XL U14123 ( .A0(\xArray[13][17] ), .A1(n8181), .B0(\xArray[1][17] ), 
        .B1(n8177), .C0(n2164), .Y(n2163) );
  OAI22XL U14124 ( .A0(n8173), .A1(n9260), .B0(n8172), .B1(n9258), .Y(n2164)
         );
  AOI221XL U14125 ( .A0(\xArray[13][18] ), .A1(n8181), .B0(\xArray[1][18] ), 
        .B1(n8177), .C0(n2155), .Y(n2154) );
  OAI22XL U14126 ( .A0(n8173), .A1(n9252), .B0(n8172), .B1(n9250), .Y(n2155)
         );
  AOI221XL U14127 ( .A0(\xArray[13][19] ), .A1(n8181), .B0(\xArray[1][19] ), 
        .B1(n8177), .C0(n2146), .Y(n2145) );
  OAI22XL U14128 ( .A0(n8173), .A1(n9244), .B0(n8172), .B1(n9242), .Y(n2146)
         );
  OAI221X1 U14129 ( .A0(\xArray[7][25] ), .A1(n8297), .B0(\xArray[11][25] ), 
        .B1(n8243), .C0(n1169), .Y(n573) );
  OAI221X1 U14130 ( .A0(\xArray[7][26] ), .A1(n8297), .B0(\xArray[11][26] ), 
        .B1(n8243), .C0(n1164), .Y(n565) );
  AOI2BB2X1 U14131 ( .B0(n9184), .B1(n8209), .A0N(\xArray[15][26] ), .A1N(
        n8256), .Y(n1164) );
  OAI221X1 U14132 ( .A0(\xArray[4][26] ), .A1(n8287), .B0(\xArray[8][26] ), 
        .B1(n8233), .C0(n2089), .Y(n1444) );
  OAI221X1 U14133 ( .A0(\xArray[4][27] ), .A1(n8287), .B0(\xArray[8][27] ), 
        .B1(n8233), .C0(n2080), .Y(n1440) );
  OAI221X1 U14134 ( .A0(\xArray[8][25] ), .A1(n8297), .B0(\xArray[12][25] ), 
        .B1(n8243), .C0(n1168), .Y(n575) );
  OAI221X1 U14135 ( .A0(\xArray[6][25] ), .A1(n8293), .B0(\xArray[10][25] ), 
        .B1(n8239), .C0(n1451), .Y(n899) );
  OA22X1 U14136 ( .A0(\xArray[14][25] ), .A1(n8271), .B0(\xArray[2][25] ), 
        .B1(n8185), .Y(n1451) );
  OAI221X1 U14137 ( .A0(\xArray[3][25] ), .A1(n8287), .B0(\xArray[7][25] ), 
        .B1(n8233), .C0(n2097), .Y(n1450) );
  OAI221X1 U14138 ( .A0(\xArray[6][26] ), .A1(n8293), .B0(\xArray[10][26] ), 
        .B1(n8239), .C0(n1447), .Y(n896) );
  OA22X1 U14139 ( .A0(\xArray[14][26] ), .A1(n8271), .B0(\xArray[2][26] ), 
        .B1(n8185), .Y(n1447) );
  OAI221X1 U14140 ( .A0(\xArray[3][26] ), .A1(n8287), .B0(\xArray[7][26] ), 
        .B1(n8233), .C0(n2088), .Y(n1446) );
  OAI221X1 U14141 ( .A0(\xArray[5][26] ), .A1(n8282), .B0(\xArray[9][26] ), 
        .B1(n8228), .C0(n1665), .Y(n1162) );
  OAI221X1 U14142 ( .A0(\xArray[5][27] ), .A1(n8282), .B0(\xArray[9][27] ), 
        .B1(n8228), .C0(n1662), .Y(n1157) );
  OAI221XL U14143 ( .A0(\xArray[9][24] ), .A1(n8291), .B0(\xArray[13][24] ), 
        .B1(n8237), .C0(n903), .Y(n582) );
  OAI221XL U14144 ( .A0(\xArray[9][25] ), .A1(n8291), .B0(\xArray[13][25] ), 
        .B1(n8237), .C0(n900), .Y(n574) );
  OAI221XL U14145 ( .A0(\xArray[2][23] ), .A1(n8287), .B0(\xArray[6][23] ), 
        .B1(n8233), .C0(n2113), .Y(n1673) );
  OAI222XL U14146 ( .A0(n653), .A1(n8339), .B0(n654), .B1(n8307), .C0(n655), 
        .C1(n7713), .Y(n648) );
  AOI221XL U14147 ( .A0(\xArray[14][15] ), .A1(n6573), .B0(\xArray[2][15] ), 
        .B1(n8361), .C0(n650), .Y(n649) );
  OAI22XL U14148 ( .A0(n8359), .A1(n9275), .B0(n6597), .B1(n9277), .Y(n650) );
  OAI222XL U14149 ( .A0(n661), .A1(n8339), .B0(n662), .B1(n8307), .C0(n663), 
        .C1(n7713), .Y(n656) );
  AOI221XL U14150 ( .A0(\xArray[14][14] ), .A1(n6573), .B0(\xArray[2][14] ), 
        .B1(n8361), .C0(n658), .Y(n657) );
  OAI22XL U14151 ( .A0(n8359), .A1(n9283), .B0(n6597), .B1(n9285), .Y(n658) );
  OAI222XL U14152 ( .A0(n669), .A1(n8339), .B0(n670), .B1(n8307), .C0(n671), 
        .C1(n7713), .Y(n664) );
  AOI221XL U14153 ( .A0(\xArray[14][13] ), .A1(n6573), .B0(\xArray[2][13] ), 
        .B1(n8361), .C0(n666), .Y(n665) );
  OAI22XL U14154 ( .A0(n8359), .A1(n9291), .B0(n8353), .B1(n9293), .Y(n666) );
  AOI221XL U14155 ( .A0(n7948), .A1(n7397), .B0(n7945), .B1(\xArray[2][11] ), 
        .C0(n4629), .Y(n4625) );
  OAI222XL U14156 ( .A0(n9306), .A1(n7943), .B0(n8708), .B1(n7938), .C0(n7935), 
        .C1(n9305), .Y(n4629) );
  OAI221XL U14157 ( .A0(n7392), .A1(n8064), .B0(n7555), .B1(n8062), .C0(n3209), 
        .Y(N28265) );
  OAI221XL U14158 ( .A0(n7392), .A1(n8141), .B0(n7555), .B1(n8139), .C0(n2710), 
        .Y(N28649) );
  OAI221XL U14159 ( .A0(n7394), .A1(n8064), .B0(n7554), .B1(n8062), .C0(n3208), 
        .Y(N28266) );
  OAI221XL U14160 ( .A0(n7394), .A1(n8141), .B0(n7554), .B1(n8139), .C0(n2708), 
        .Y(N28650) );
  OAI221XL U14161 ( .A0(n7396), .A1(n8064), .B0(n7553), .B1(n8062), .C0(n3207), 
        .Y(N28267) );
  OAI221XL U14162 ( .A0(n7396), .A1(n8141), .B0(n7553), .B1(n8139), .C0(n2706), 
        .Y(N28651) );
  OAI221XL U14163 ( .A0(n7398), .A1(n8064), .B0(n7552), .B1(n8062), .C0(n3206), 
        .Y(N28268) );
  OAI221XL U14164 ( .A0(n7398), .A1(n8141), .B0(n7552), .B1(n8139), .C0(n2704), 
        .Y(N28652) );
  MX4X1 U14165 ( .A(n6808), .B(n6806), .C(n6807), .D(n6805), .S0(n7005), .S1(
        n7003), .Y(N25579) );
  MX4X1 U14166 ( .A(n6804), .B(n6802), .C(n6803), .D(n6801), .S0(n7005), .S1(
        n7003), .Y(N25580) );
  AND4X1 U14167 ( .A(n4677), .B(n4678), .C(n4679), .D(n4680), .Y(n2496) );
  AOI221XL U14168 ( .A0(n7962), .A1(\xArray[9][8] ), .B0(\xArray[8][8] ), .B1(
        n7960), .C0(n4681), .Y(n4680) );
  AOI221XL U14169 ( .A0(n7949), .A1(n7391), .B0(n7944), .B1(\xArray[2][8] ), 
        .C0(n4683), .Y(n4679) );
  AND4X1 U14170 ( .A(n4659), .B(n4660), .C(n4661), .D(n4662), .Y(n2493) );
  AOI221XL U14171 ( .A0(n7962), .A1(\xArray[9][9] ), .B0(\xArray[8][9] ), .B1(
        n3660), .C0(n4663), .Y(n4662) );
  AOI221XL U14172 ( .A0(n7947), .A1(n7393), .B0(n7946), .B1(\xArray[2][9] ), 
        .C0(n4665), .Y(n4661) );
  AND4X1 U14173 ( .A(n4641), .B(n4642), .C(n4643), .D(n4644), .Y(n2490) );
  AOI221XL U14174 ( .A0(n7962), .A1(\xArray[9][10] ), .B0(\xArray[8][10] ), 
        .B1(n3660), .C0(n4645), .Y(n4644) );
  AOI221XL U14175 ( .A0(n7949), .A1(n7395), .B0(n7945), .B1(\xArray[2][10] ), 
        .C0(n4647), .Y(n4643) );
  AND4X1 U14176 ( .A(n4623), .B(n4624), .C(n4625), .D(n4626), .Y(n2487) );
  AOI221XL U14177 ( .A0(n7962), .A1(\xArray[9][11] ), .B0(\xArray[8][11] ), 
        .B1(n3660), .C0(n4627), .Y(n4626) );
  AOI221XL U14178 ( .A0(n8711), .A1(n7992), .B0(n8712), .B1(n8029), .C0(n4632), 
        .Y(n4624) );
  MX4X1 U14179 ( .A(\bArray[12][22] ), .B(\bArray[13][22] ), .C(
        \bArray[14][22] ), .D(\bArray[15][22] ), .S0(n7207), .S1(n7219), .Y(
        n7032) );
  MX4X1 U14180 ( .A(\bArray[8][22] ), .B(\bArray[9][22] ), .C(\bArray[10][22] ), .D(\bArray[11][22] ), .S0(n7207), .S1(n7219), .Y(n7033) );
  MX4X1 U14181 ( .A(\bArray[4][22] ), .B(\bArray[5][22] ), .C(\bArray[6][22] ), 
        .D(\bArray[7][22] ), .S0(n7207), .S1(n7219), .Y(n7034) );
  OAI221X1 U14182 ( .A0(\xArray[7][27] ), .A1(n8298), .B0(\xArray[11][27] ), 
        .B1(n8232), .C0(n1159), .Y(n557) );
  AOI2BB2X1 U14183 ( .B0(n9176), .B1(n8209), .A0N(\xArray[15][27] ), .A1N(
        n8256), .Y(n1159) );
  OAI221X1 U14184 ( .A0(\xArray[7][28] ), .A1(n8298), .B0(\xArray[11][28] ), 
        .B1(n8232), .C0(n1154), .Y(n549) );
  OAI221X1 U14185 ( .A0(\xArray[4][28] ), .A1(n8287), .B0(\xArray[8][28] ), 
        .B1(n8233), .C0(n2071), .Y(n1436) );
  OAI221X1 U14186 ( .A0(\xArray[4][29] ), .A1(n8288), .B0(\xArray[8][29] ), 
        .B1(n8234), .C0(n2062), .Y(n1432) );
  OA22X1 U14187 ( .A0(\xArray[0][29] ), .A1(n8192), .B0(\xArray[12][29] ), 
        .B1(n8266), .Y(n2062) );
  OAI221X1 U14188 ( .A0(\xArray[8][26] ), .A1(n8298), .B0(\xArray[12][26] ), 
        .B1(n8236), .C0(n1163), .Y(n567) );
  OA22X1 U14189 ( .A0(\xArray[4][26] ), .A1(n8197), .B0(\xArray[0][26] ), .B1(
        n8267), .Y(n1163) );
  OAI221X1 U14190 ( .A0(\xArray[8][27] ), .A1(n8298), .B0(\xArray[12][27] ), 
        .B1(n8236), .C0(n1158), .Y(n559) );
  OA22X1 U14191 ( .A0(\xArray[4][27] ), .A1(n8197), .B0(\xArray[0][27] ), .B1(
        n8267), .Y(n1158) );
  OAI221X1 U14192 ( .A0(\xArray[3][27] ), .A1(n8287), .B0(\xArray[7][27] ), 
        .B1(n8233), .C0(n2079), .Y(n1442) );
  OAI221X1 U14193 ( .A0(\xArray[5][28] ), .A1(n8282), .B0(\xArray[9][28] ), 
        .B1(n8228), .C0(n1659), .Y(n1152) );
  OA22X1 U14194 ( .A0(\xArray[1][28] ), .A1(n8188), .B0(\xArray[13][28] ), 
        .B1(n8262), .Y(n1659) );
  OAI221X1 U14195 ( .A0(\xArray[5][29] ), .A1(n8282), .B0(\xArray[9][29] ), 
        .B1(n8228), .C0(n1656), .Y(n1147) );
  OA22X1 U14196 ( .A0(\xArray[1][29] ), .A1(n8188), .B0(\xArray[13][29] ), 
        .B1(n8262), .Y(n1656) );
  OAI221XL U14197 ( .A0(\xArray[2][24] ), .A1(n8287), .B0(\xArray[6][24] ), 
        .B1(n8233), .C0(n2104), .Y(n1670) );
  OAI221XL U14198 ( .A0(\xArray[2][25] ), .A1(n8287), .B0(\xArray[6][25] ), 
        .B1(n8233), .C0(n2095), .Y(n1667) );
  OAI221XL U14199 ( .A0(\xArray[2][26] ), .A1(n8287), .B0(\xArray[6][26] ), 
        .B1(n8233), .C0(n2086), .Y(n1664) );
  OAI222XL U14200 ( .A0(n645), .A1(n8339), .B0(n646), .B1(n8307), .C0(n647), 
        .C1(n7713), .Y(n640) );
  AOI221XL U14201 ( .A0(\xArray[14][16] ), .A1(n6573), .B0(\xArray[2][16] ), 
        .B1(n8360), .C0(n642), .Y(n641) );
  OAI22XL U14202 ( .A0(n8359), .A1(n9267), .B0(n6597), .B1(n9269), .Y(n642) );
  OAI221XL U14203 ( .A0(n7380), .A1(n8064), .B0(n7561), .B1(n8062), .C0(n3215), 
        .Y(N28259) );
  OAI221XL U14204 ( .A0(n7380), .A1(n8141), .B0(n7561), .B1(n8139), .C0(n2722), 
        .Y(N28643) );
  OAI221XL U14205 ( .A0(n7382), .A1(n8064), .B0(n7560), .B1(n8062), .C0(n3214), 
        .Y(N28260) );
  OAI221XL U14206 ( .A0(n7382), .A1(n8141), .B0(n7560), .B1(n8139), .C0(n2720), 
        .Y(N28644) );
  OAI221XL U14207 ( .A0(n7384), .A1(n8064), .B0(n7559), .B1(n8062), .C0(n3213), 
        .Y(N28261) );
  OAI221XL U14208 ( .A0(n7384), .A1(n8141), .B0(n7559), .B1(n8139), .C0(n2718), 
        .Y(N28645) );
  OAI221XL U14209 ( .A0(n7386), .A1(n8064), .B0(n7558), .B1(n8062), .C0(n3212), 
        .Y(N28262) );
  OAI221XL U14210 ( .A0(n7386), .A1(n8141), .B0(n7558), .B1(n8139), .C0(n2716), 
        .Y(N28646) );
  OAI221XL U14211 ( .A0(n7388), .A1(n8064), .B0(n7557), .B1(n8062), .C0(n3211), 
        .Y(N28263) );
  OAI221XL U14212 ( .A0(n7388), .A1(n8141), .B0(n7557), .B1(n8139), .C0(n2714), 
        .Y(N28647) );
  OAI221XL U14213 ( .A0(n7390), .A1(n8064), .B0(n7556), .B1(n8062), .C0(n3210), 
        .Y(N28264) );
  OAI221XL U14214 ( .A0(n7390), .A1(n8141), .B0(n7556), .B1(n8139), .C0(n2712), 
        .Y(N28648) );
  MX4X1 U14215 ( .A(n6816), .B(n6814), .C(n6815), .D(n6813), .S0(n7005), .S1(
        n7003), .Y(N25577) );
  MX4X1 U14216 ( .A(n6812), .B(n6810), .C(n6811), .D(n6809), .S0(n7005), .S1(
        n7003), .Y(N25578) );
  AND4X1 U14217 ( .A(n4785), .B(n4786), .C(n4787), .D(n4788), .Y(n2514) );
  AOI221XL U14218 ( .A0(n7963), .A1(\xArray[9][2] ), .B0(\xArray[8][2] ), .B1(
        n7959), .C0(n4789), .Y(n4788) );
  AOI221XL U14219 ( .A0(n7948), .A1(n7379), .B0(n3667), .B1(\xArray[2][2] ), 
        .C0(n4791), .Y(n4787) );
  AND4X1 U14220 ( .A(n4767), .B(n4768), .C(n4769), .D(n4770), .Y(n2511) );
  AOI221XL U14221 ( .A0(n7963), .A1(\xArray[9][3] ), .B0(\xArray[8][3] ), .B1(
        n7959), .C0(n4771), .Y(n4770) );
  AOI221XL U14222 ( .A0(n7949), .A1(n7381), .B0(n7946), .B1(\xArray[2][3] ), 
        .C0(n4773), .Y(n4769) );
  AND4X1 U14223 ( .A(n4749), .B(n4750), .C(n4751), .D(n4752), .Y(n2508) );
  AOI221XL U14224 ( .A0(n3659), .A1(\xArray[9][4] ), .B0(\xArray[8][4] ), .B1(
        n7959), .C0(n4753), .Y(n4752) );
  AOI221XL U14225 ( .A0(n7947), .A1(n7383), .B0(n7944), .B1(\xArray[2][4] ), 
        .C0(n4755), .Y(n4751) );
  AND4X1 U14226 ( .A(n4731), .B(n4732), .C(n4733), .D(n4734), .Y(n2505) );
  AOI221XL U14227 ( .A0(n3659), .A1(\xArray[9][5] ), .B0(\xArray[8][5] ), .B1(
        n7959), .C0(n4735), .Y(n4734) );
  AOI221XL U14228 ( .A0(n7949), .A1(n7385), .B0(n7944), .B1(\xArray[2][5] ), 
        .C0(n4737), .Y(n4733) );
  AND4X1 U14229 ( .A(n4713), .B(n4714), .C(n4715), .D(n4716), .Y(n2502) );
  AOI221XL U14230 ( .A0(n3659), .A1(\xArray[9][6] ), .B0(\xArray[8][6] ), .B1(
        n7959), .C0(n4717), .Y(n4716) );
  AOI221XL U14231 ( .A0(n7948), .A1(n7387), .B0(n7945), .B1(\xArray[2][6] ), 
        .C0(n4719), .Y(n4715) );
  AND4X1 U14232 ( .A(n4695), .B(n4696), .C(n4697), .D(n4698), .Y(n2499) );
  AOI221XL U14233 ( .A0(n7964), .A1(\xArray[9][7] ), .B0(\xArray[8][7] ), .B1(
        n7960), .C0(n4699), .Y(n4698) );
  AOI221XL U14234 ( .A0(n7948), .A1(n7389), .B0(n7944), .B1(\xArray[2][7] ), 
        .C0(n4701), .Y(n4697) );
  OAI221X1 U14235 ( .A0(\xArray[6][27] ), .A1(n8293), .B0(\xArray[10][27] ), 
        .B1(n8239), .C0(n1443), .Y(n893) );
  OAI221X1 U14236 ( .A0(\xArray[6][28] ), .A1(n8294), .B0(\xArray[10][28] ), 
        .B1(n8240), .C0(n1439), .Y(n890) );
  OA22X1 U14237 ( .A0(\xArray[14][28] ), .A1(n8271), .B0(\xArray[2][28] ), 
        .B1(n8185), .Y(n1439) );
  OAI221XL U14238 ( .A0(\xArray[9][26] ), .A1(n8291), .B0(\xArray[13][26] ), 
        .B1(n8237), .C0(n897), .Y(n566) );
  OAI221XL U14239 ( .A0(\xArray[9][27] ), .A1(n8291), .B0(\xArray[13][27] ), 
        .B1(n8237), .C0(n894), .Y(n558) );
  OAI221X1 U14240 ( .A0(\xArray[3][28] ), .A1(n8287), .B0(\xArray[7][28] ), 
        .B1(n8233), .C0(n2070), .Y(n1438) );
  AOI221XL U14241 ( .A0(\xArray[13][20] ), .A1(n8181), .B0(\xArray[1][20] ), 
        .B1(n8177), .C0(n2137), .Y(n2136) );
  OAI22XL U14242 ( .A0(n1749), .A1(n9236), .B0(n8172), .B1(n9234), .Y(n2137)
         );
  AOI221XL U14243 ( .A0(\xArray[13][21] ), .A1(n8181), .B0(\xArray[1][21] ), 
        .B1(n8177), .C0(n2128), .Y(n2127) );
  OAI22XL U14244 ( .A0(n8173), .A1(n9228), .B0(n8172), .B1(n9226), .Y(n2128)
         );
  AOI221XL U14245 ( .A0(\xArray[13][22] ), .A1(n8181), .B0(\xArray[1][22] ), 
        .B1(n8177), .C0(n2119), .Y(n2118) );
  OA22X1 U14246 ( .A0(n8312), .A1(n1462), .B0(n7729), .B1(n1676), .Y(n2117) );
  OAI22XL U14247 ( .A0(n8173), .A1(n9220), .B0(n8172), .B1(n9218), .Y(n2119)
         );
  AOI221XL U14248 ( .A0(\xArray[13][23] ), .A1(n8181), .B0(\xArray[1][23] ), 
        .B1(n8177), .C0(n2110), .Y(n2109) );
  OA22X1 U14249 ( .A0(n8312), .A1(n1458), .B0(n7729), .B1(n1673), .Y(n2108) );
  OAI22XL U14250 ( .A0(n8173), .A1(n9212), .B0(n8172), .B1(n9210), .Y(n2110)
         );
  OAI221X1 U14251 ( .A0(\xArray[7][29] ), .A1(n8298), .B0(\xArray[11][29] ), 
        .B1(n8232), .C0(n1149), .Y(n541) );
  OAI221X1 U14252 ( .A0(\xArray[7][30] ), .A1(n8298), .B0(\xArray[11][30] ), 
        .B1(n8224), .C0(n1144), .Y(n533) );
  OAI221X1 U14253 ( .A0(\xArray[4][30] ), .A1(n8288), .B0(\xArray[8][30] ), 
        .B1(n8234), .C0(n2053), .Y(n1428) );
  OAI221X1 U14254 ( .A0(\xArray[8][28] ), .A1(n8298), .B0(\xArray[12][28] ), 
        .B1(n8241), .C0(n1153), .Y(n551) );
  OAI221X1 U14255 ( .A0(\xArray[8][29] ), .A1(n8298), .B0(\xArray[12][29] ), 
        .B1(n8224), .C0(n1148), .Y(n543) );
  OAI221X1 U14256 ( .A0(\xArray[5][30] ), .A1(n8282), .B0(\xArray[9][30] ), 
        .B1(n8228), .C0(n1653), .Y(n1142) );
  OAI221XL U14257 ( .A0(\xArray[2][27] ), .A1(n8287), .B0(\xArray[6][27] ), 
        .B1(n8233), .C0(n2077), .Y(n1661) );
  OAI221XL U14258 ( .A0(\xArray[2][28] ), .A1(n8288), .B0(\xArray[6][28] ), 
        .B1(n8234), .C0(n2068), .Y(n1658) );
  AOI2BB2X1 U14259 ( .B0(n9174), .B1(n8208), .A0N(\xArray[10][28] ), .A1N(
        n8256), .Y(n2068) );
  OAI222XL U14260 ( .A0(n621), .A1(n8339), .B0(n622), .B1(n8307), .C0(n623), 
        .C1(n7713), .Y(n616) );
  AOI221XL U14261 ( .A0(\xArray[14][19] ), .A1(n6573), .B0(\xArray[2][19] ), 
        .B1(n8360), .C0(n618), .Y(n617) );
  OAI22XL U14262 ( .A0(n8359), .A1(n9243), .B0(n6597), .B1(n9245), .Y(n618) );
  OAI222XL U14263 ( .A0(n629), .A1(n8339), .B0(n630), .B1(n8307), .C0(n631), 
        .C1(n7713), .Y(n624) );
  AOI221XL U14264 ( .A0(\xArray[14][18] ), .A1(n6573), .B0(\xArray[2][18] ), 
        .B1(n8360), .C0(n626), .Y(n625) );
  OAI22XL U14265 ( .A0(n8359), .A1(n9251), .B0(n6597), .B1(n9253), .Y(n626) );
  OAI222XL U14266 ( .A0(n637), .A1(n8339), .B0(n638), .B1(n8307), .C0(n639), 
        .C1(n7713), .Y(n632) );
  AOI221XL U14267 ( .A0(\xArray[14][17] ), .A1(n6573), .B0(\xArray[2][17] ), 
        .B1(n8360), .C0(n634), .Y(n633) );
  OAI22XL U14268 ( .A0(n8359), .A1(n9259), .B0(n6597), .B1(n9261), .Y(n634) );
  AOI221XL U14269 ( .A0(n7947), .A1(n7375), .B0(n7944), .B1(\xArray[2][0] ), 
        .C0(n4847), .Y(n4836) );
  OAI222XL U14270 ( .A0(n9394), .A1(n3669), .B0(n8763), .B1(n7938), .C0(n7935), 
        .C1(n9393), .Y(n4847) );
  AOI221XL U14271 ( .A0(n7947), .A1(n7377), .B0(n7945), .B1(\xArray[2][1] ), 
        .C0(n4809), .Y(n4805) );
  OAI222XL U14272 ( .A0(n9386), .A1(n7943), .B0(n8758), .B1(n7939), .C0(n7935), 
        .C1(n9385), .Y(n4809) );
  OAI221XL U14273 ( .A0(n7376), .A1(n8064), .B0(n7563), .B1(n8062), .C0(n3217), 
        .Y(N28257) );
  OAI221XL U14274 ( .A0(n7376), .A1(n8141), .B0(n7563), .B1(n8139), .C0(n2726), 
        .Y(N28641) );
  OAI221XL U14275 ( .A0(n7378), .A1(n8064), .B0(n7562), .B1(n8062), .C0(n3216), 
        .Y(N28258) );
  OAI221XL U14276 ( .A0(n7378), .A1(n8141), .B0(n7562), .B1(n8139), .C0(n2724), 
        .Y(N28642) );
  MX4X1 U14277 ( .A(n6824), .B(n6822), .C(n6823), .D(n6821), .S0(n7005), .S1(
        n7003), .Y(N25575) );
  MX4X1 U14278 ( .A(n6820), .B(n6818), .C(n6819), .D(n6817), .S0(n7005), .S1(
        n7003), .Y(N25576) );
  AND4X1 U14279 ( .A(n4834), .B(n4835), .C(n4836), .D(n4837), .Y(n2520) );
  AOI221XL U14280 ( .A0(n7963), .A1(\xArray[9][0] ), .B0(\xArray[8][0] ), .B1(
        n7959), .C0(n4838), .Y(n4837) );
  AOI221XL U14281 ( .A0(n8766), .A1(n7994), .B0(n8767), .B1(n8031), .C0(n4857), 
        .Y(n4835) );
  AND4X1 U14282 ( .A(n4803), .B(n4804), .C(n4805), .D(n4806), .Y(n2517) );
  AOI221XL U14283 ( .A0(n7963), .A1(\xArray[9][1] ), .B0(\xArray[8][1] ), .B1(
        n7961), .C0(n4807), .Y(n4806) );
  AOI221XL U14284 ( .A0(n8761), .A1(n7992), .B0(n8762), .B1(n8029), .C0(n4812), 
        .Y(n4804) );
  OAI221X1 U14285 ( .A0(\xArray[6][29] ), .A1(n8294), .B0(\xArray[10][29] ), 
        .B1(n8240), .C0(n1435), .Y(n887) );
  OA22X1 U14286 ( .A0(\xArray[14][29] ), .A1(n8271), .B0(\xArray[2][29] ), 
        .B1(n8185), .Y(n1435) );
  OAI221X1 U14287 ( .A0(\xArray[6][30] ), .A1(n8294), .B0(\xArray[10][30] ), 
        .B1(n8240), .C0(n1431), .Y(n884) );
  OAI221XL U14288 ( .A0(\xArray[9][28] ), .A1(n8291), .B0(\xArray[13][28] ), 
        .B1(n8237), .C0(n891), .Y(n550) );
  OAI221XL U14289 ( .A0(\xArray[9][29] ), .A1(n8291), .B0(\xArray[13][29] ), 
        .B1(n8237), .C0(n888), .Y(n542) );
  OAI221X1 U14290 ( .A0(\xArray[3][29] ), .A1(n8288), .B0(\xArray[7][29] ), 
        .B1(n8234), .C0(n2061), .Y(n1434) );
  OA22X1 U14291 ( .A0(\xArray[15][29] ), .A1(n8192), .B0(\xArray[11][29] ), 
        .B1(n8266), .Y(n2061) );
  OAI221X1 U14292 ( .A0(\xArray[3][30] ), .A1(n8288), .B0(\xArray[7][30] ), 
        .B1(n8234), .C0(n2052), .Y(n1430) );
  MX4X1 U14293 ( .A(\bArray[12][25] ), .B(\bArray[13][25] ), .C(
        \bArray[14][25] ), .D(\bArray[15][25] ), .S0(n7208), .S1(n7220), .Y(
        n7044) );
  MX4X1 U14294 ( .A(\bArray[8][25] ), .B(\bArray[9][25] ), .C(\bArray[10][25] ), .D(\bArray[11][25] ), .S0(n7208), .S1(n7220), .Y(n7045) );
  MX4X1 U14295 ( .A(\bArray[4][25] ), .B(\bArray[5][25] ), .C(\bArray[6][25] ), 
        .D(\bArray[7][25] ), .S0(n7208), .S1(n7220), .Y(n7046) );
  OAI221X1 U14296 ( .A0(\xArray[7][31] ), .A1(n8298), .B0(\xArray[11][31] ), 
        .B1(n8232), .C0(n1139), .Y(n525) );
  OAI221X1 U14297 ( .A0(\xArray[4][31] ), .A1(n8288), .B0(\xArray[8][31] ), 
        .B1(n8234), .C0(n2044), .Y(n1424) );
  OAI221X1 U14298 ( .A0(\xArray[4][32] ), .A1(n8288), .B0(\xArray[8][32] ), 
        .B1(n8234), .C0(n2035), .Y(n1420) );
  OAI221X1 U14299 ( .A0(\xArray[8][30] ), .A1(n8298), .B0(\xArray[12][30] ), 
        .B1(n8232), .C0(n1143), .Y(n535) );
  OAI221X1 U14300 ( .A0(\xArray[8][31] ), .A1(n8289), .B0(\xArray[12][31] ), 
        .B1(n8235), .C0(n1138), .Y(n527) );
  OA22X1 U14301 ( .A0(\xArray[4][31] ), .A1(n8197), .B0(\xArray[0][31] ), .B1(
        n8267), .Y(n1138) );
  OAI221X1 U14302 ( .A0(\xArray[6][31] ), .A1(n8294), .B0(\xArray[10][31] ), 
        .B1(n8240), .C0(n1427), .Y(n881) );
  OAI221X1 U14303 ( .A0(\xArray[6][32] ), .A1(n8294), .B0(\xArray[10][32] ), 
        .B1(n8240), .C0(n1423), .Y(n878) );
  OAI221X1 U14304 ( .A0(\xArray[5][31] ), .A1(n8282), .B0(\xArray[9][31] ), 
        .B1(n8228), .C0(n1650), .Y(n1137) );
  OAI221X1 U14305 ( .A0(\xArray[5][32] ), .A1(n8282), .B0(\xArray[9][32] ), 
        .B1(n8228), .C0(n1647), .Y(n1132) );
  OA22X1 U14306 ( .A0(\xArray[1][32] ), .A1(n8200), .B0(\xArray[13][32] ), 
        .B1(n8260), .Y(n1647) );
  OAI221XL U14307 ( .A0(\xArray[2][29] ), .A1(n8288), .B0(\xArray[6][29] ), 
        .B1(n8234), .C0(n2059), .Y(n1655) );
  OAI221XL U14308 ( .A0(\xArray[2][30] ), .A1(n8288), .B0(\xArray[6][30] ), 
        .B1(n8234), .C0(n2050), .Y(n1652) );
  OAI222XL U14309 ( .A0(n613), .A1(n8339), .B0(n614), .B1(n8307), .C0(n615), 
        .C1(n7713), .Y(n608) );
  AOI221XL U14310 ( .A0(\xArray[14][20] ), .A1(n6573), .B0(\xArray[2][20] ), 
        .B1(n8360), .C0(n610), .Y(n609) );
  OAI22XL U14311 ( .A0(n8359), .A1(n9235), .B0(n6597), .B1(n9237), .Y(n610) );
  MX4X1 U14312 ( .A(n6832), .B(n6830), .C(n6831), .D(n6829), .S0(n8411), .S1(
        n7004), .Y(N25573) );
  MX4X1 U14313 ( .A(n6828), .B(n6826), .C(n6827), .D(n6825), .S0(n8411), .S1(
        n8412), .Y(N25574) );
  MX4X1 U14314 ( .A(\bArray[0][25] ), .B(\bArray[1][25] ), .C(\bArray[2][25] ), 
        .D(\bArray[3][25] ), .S0(n7208), .S1(n7220), .Y(n7047) );
  OAI221XL U14315 ( .A0(\xArray[9][30] ), .A1(n8291), .B0(\xArray[13][30] ), 
        .B1(n8237), .C0(n885), .Y(n534) );
  OAI221XL U14316 ( .A0(\xArray[9][31] ), .A1(n8291), .B0(\xArray[13][31] ), 
        .B1(n8237), .C0(n882), .Y(n526) );
  OAI221X1 U14317 ( .A0(\xArray[3][31] ), .A1(n8288), .B0(\xArray[7][31] ), 
        .B1(n8234), .C0(n2043), .Y(n1426) );
  OAI221X1 U14318 ( .A0(\xArray[3][32] ), .A1(n8288), .B0(\xArray[7][32] ), 
        .B1(n8234), .C0(n2034), .Y(n1422) );
  AOI221XL U14319 ( .A0(\xArray[13][24] ), .A1(n8181), .B0(\xArray[1][24] ), 
        .B1(n8177), .C0(n2101), .Y(n2100) );
  OA22X1 U14320 ( .A0(n8312), .A1(n1454), .B0(n7729), .B1(n1670), .Y(n2099) );
  OAI22XL U14321 ( .A0(n8173), .A1(n9204), .B0(n8172), .B1(n9202), .Y(n2101)
         );
  AOI221XL U14322 ( .A0(\xArray[13][25] ), .A1(n8181), .B0(\xArray[1][25] ), 
        .B1(n8177), .C0(n2092), .Y(n2091) );
  OA22X1 U14323 ( .A0(n8312), .A1(n1450), .B0(n7729), .B1(n1667), .Y(n2090) );
  OAI22XL U14324 ( .A0(n8173), .A1(n9196), .B0(n8172), .B1(n9194), .Y(n2092)
         );
  AOI221XL U14325 ( .A0(\xArray[13][26] ), .A1(n8181), .B0(\xArray[1][26] ), 
        .B1(n8177), .C0(n2083), .Y(n2082) );
  OA22X1 U14326 ( .A0(n8312), .A1(n1446), .B0(n7729), .B1(n1664), .Y(n2081) );
  OAI22XL U14327 ( .A0(n8173), .A1(n9188), .B0(n8170), .B1(n9186), .Y(n2083)
         );
  AOI221XL U14328 ( .A0(\xArray[13][27] ), .A1(n8181), .B0(\xArray[1][27] ), 
        .B1(n8177), .C0(n2074), .Y(n2073) );
  OA22X1 U14329 ( .A0(n8312), .A1(n1442), .B0(n7729), .B1(n1661), .Y(n2072) );
  OAI22XL U14330 ( .A0(n8174), .A1(n9180), .B0(n8172), .B1(n9178), .Y(n2074)
         );
  OAI221X1 U14331 ( .A0(\xArray[7][32] ), .A1(n8290), .B0(\xArray[11][32] ), 
        .B1(n8225), .C0(n1134), .Y(n517) );
  AOI2BB2X1 U14332 ( .B0(n9136), .B1(n8212), .A0N(\xArray[15][32] ), .A1N(
        n8256), .Y(n1134) );
  OAI221X1 U14333 ( .A0(\xArray[7][33] ), .A1(n8290), .B0(\xArray[11][33] ), 
        .B1(n8225), .C0(n1129), .Y(n509) );
  OAI221X1 U14334 ( .A0(\xArray[7][34] ), .A1(n8290), .B0(\xArray[11][34] ), 
        .B1(n8226), .C0(n1124), .Y(n501) );
  OAI221X1 U14335 ( .A0(\xArray[4][33] ), .A1(n8288), .B0(\xArray[8][33] ), 
        .B1(n8234), .C0(n2026), .Y(n1416) );
  OAI221X1 U14336 ( .A0(\xArray[4][34] ), .A1(n8288), .B0(\xArray[8][34] ), 
        .B1(n8234), .C0(n2017), .Y(n1412) );
  OAI221X1 U14337 ( .A0(\xArray[8][32] ), .A1(n8286), .B0(\xArray[12][32] ), 
        .B1(n8230), .C0(n1133), .Y(n519) );
  OA22X1 U14338 ( .A0(\xArray[4][32] ), .A1(n8197), .B0(\xArray[0][32] ), .B1(
        n8267), .Y(n1133) );
  OAI221X1 U14339 ( .A0(\xArray[8][33] ), .A1(n8292), .B0(\xArray[12][33] ), 
        .B1(n8230), .C0(n1128), .Y(n511) );
  OAI221X1 U14340 ( .A0(\xArray[6][33] ), .A1(n8294), .B0(\xArray[10][33] ), 
        .B1(n8240), .C0(n1419), .Y(n875) );
  OAI221X1 U14341 ( .A0(\xArray[6][34] ), .A1(n8294), .B0(\xArray[10][34] ), 
        .B1(n8240), .C0(n1415), .Y(n872) );
  OAI221X1 U14342 ( .A0(\xArray[5][33] ), .A1(n8282), .B0(\xArray[9][33] ), 
        .B1(n8228), .C0(n1644), .Y(n1127) );
  OA22X1 U14343 ( .A0(\xArray[1][33] ), .A1(n8200), .B0(\xArray[13][33] ), 
        .B1(n8257), .Y(n1644) );
  OAI221X1 U14344 ( .A0(\xArray[5][34] ), .A1(n8282), .B0(\xArray[9][34] ), 
        .B1(n8228), .C0(n1641), .Y(n1122) );
  OA22X1 U14345 ( .A0(\xArray[1][34] ), .A1(n8200), .B0(\xArray[13][34] ), 
        .B1(n8273), .Y(n1641) );
  OAI221XL U14346 ( .A0(\xArray[9][32] ), .A1(n8291), .B0(\xArray[13][32] ), 
        .B1(n8237), .C0(n879), .Y(n518) );
  OAI221XL U14347 ( .A0(\xArray[9][33] ), .A1(n8291), .B0(\xArray[13][33] ), 
        .B1(n8237), .C0(n876), .Y(n510) );
  OAI221XL U14348 ( .A0(\xArray[2][31] ), .A1(n8288), .B0(\xArray[6][31] ), 
        .B1(n8234), .C0(n2041), .Y(n1649) );
  OAI221XL U14349 ( .A0(\xArray[2][32] ), .A1(n8288), .B0(\xArray[6][32] ), 
        .B1(n8234), .C0(n2032), .Y(n1646) );
  OAI222XL U14350 ( .A0(n589), .A1(n8339), .B0(n590), .B1(n8307), .C0(n591), 
        .C1(n7713), .Y(n584) );
  AOI221XL U14351 ( .A0(\xArray[14][23] ), .A1(n6573), .B0(\xArray[2][23] ), 
        .B1(n8360), .C0(n586), .Y(n585) );
  OAI22XL U14352 ( .A0(n8359), .A1(n9211), .B0(n6597), .B1(n9213), .Y(n586) );
  OAI222XL U14353 ( .A0(n597), .A1(n8339), .B0(n598), .B1(n8307), .C0(n599), 
        .C1(n7713), .Y(n592) );
  AOI221XL U14354 ( .A0(\xArray[14][22] ), .A1(n6573), .B0(\xArray[2][22] ), 
        .B1(n8360), .C0(n594), .Y(n593) );
  OAI22XL U14355 ( .A0(n8359), .A1(n9219), .B0(n6597), .B1(n9221), .Y(n594) );
  OAI222XL U14356 ( .A0(n605), .A1(n8339), .B0(n606), .B1(n8307), .C0(n607), 
        .C1(n7713), .Y(n600) );
  AOI221XL U14357 ( .A0(\xArray[14][21] ), .A1(n6573), .B0(\xArray[2][21] ), 
        .B1(n8360), .C0(n602), .Y(n601) );
  OAI22XL U14358 ( .A0(n8359), .A1(n9227), .B0(n6597), .B1(n9229), .Y(n602) );
  MX4X1 U14359 ( .A(n6840), .B(n6838), .C(n6839), .D(n6837), .S0(n7006), .S1(
        n7004), .Y(N25571) );
  MX4X1 U14360 ( .A(n6836), .B(n6834), .C(n6835), .D(n6833), .S0(n7006), .S1(
        n7004), .Y(N25572) );
  OAI221X1 U14361 ( .A0(\xArray[3][33] ), .A1(n8288), .B0(\xArray[7][33] ), 
        .B1(n8234), .C0(n2025), .Y(n1418) );
  OAI221X1 U14362 ( .A0(\xArray[3][34] ), .A1(n8288), .B0(\xArray[7][34] ), 
        .B1(n8234), .C0(n2016), .Y(n1414) );
  MX4X1 U14363 ( .A(\bArray[8][28] ), .B(\bArray[9][28] ), .C(\bArray[10][28] ), .D(\bArray[11][28] ), .S0(n7209), .S1(n7221), .Y(n7057) );
  MX4X1 U14364 ( .A(\bArray[4][28] ), .B(\bArray[5][28] ), .C(\bArray[6][28] ), 
        .D(\bArray[7][28] ), .S0(n7209), .S1(n7221), .Y(n7058) );
  MX4X1 U14365 ( .A(\bArray[4][31] ), .B(\bArray[5][31] ), .C(\bArray[6][31] ), 
        .D(\bArray[7][31] ), .S0(n7210), .S1(n8409), .Y(n7070) );
  OAI221X1 U14366 ( .A0(\xArray[7][35] ), .A1(n8290), .B0(\xArray[11][35] ), 
        .B1(n8226), .C0(n1119), .Y(n493) );
  OAI221X1 U14367 ( .A0(\xArray[7][36] ), .A1(n8290), .B0(\xArray[11][36] ), 
        .B1(n8226), .C0(n1114), .Y(n485) );
  OAI221X1 U14368 ( .A0(\xArray[4][35] ), .A1(n8283), .B0(\xArray[8][35] ), 
        .B1(n8235), .C0(n2008), .Y(n1408) );
  OA22X1 U14369 ( .A0(\xArray[0][35] ), .A1(n8192), .B0(\xArray[12][35] ), 
        .B1(n8265), .Y(n2008) );
  OAI221X1 U14370 ( .A0(\xArray[4][36] ), .A1(n8283), .B0(\xArray[8][36] ), 
        .B1(n8235), .C0(n1999), .Y(n1404) );
  OAI221X1 U14371 ( .A0(\xArray[4][37] ), .A1(n8280), .B0(\xArray[8][37] ), 
        .B1(n8235), .C0(n1990), .Y(n1400) );
  OAI221X1 U14372 ( .A0(\xArray[8][34] ), .A1(n8286), .B0(\xArray[12][34] ), 
        .B1(n8226), .C0(n1123), .Y(n503) );
  OAI221X1 U14373 ( .A0(\xArray[8][35] ), .A1(n8286), .B0(\xArray[12][35] ), 
        .B1(n8226), .C0(n1118), .Y(n495) );
  OAI221X1 U14374 ( .A0(\xArray[6][35] ), .A1(n8294), .B0(\xArray[10][35] ), 
        .B1(n8240), .C0(n1411), .Y(n869) );
  OAI221X1 U14375 ( .A0(\xArray[6][36] ), .A1(n8294), .B0(\xArray[10][36] ), 
        .B1(n8240), .C0(n1407), .Y(n866) );
  OAI221X1 U14376 ( .A0(\xArray[5][35] ), .A1(n8282), .B0(\xArray[9][35] ), 
        .B1(n8228), .C0(n1638), .Y(n1117) );
  OA22X1 U14377 ( .A0(\xArray[1][35] ), .A1(n8200), .B0(\xArray[13][35] ), 
        .B1(n8268), .Y(n1638) );
  OAI221X1 U14378 ( .A0(\xArray[5][36] ), .A1(n8282), .B0(\xArray[9][36] ), 
        .B1(n8228), .C0(n1635), .Y(n1112) );
  OA22X1 U14379 ( .A0(\xArray[1][36] ), .A1(n8200), .B0(\xArray[13][36] ), 
        .B1(n8257), .Y(n1635) );
  OAI221X1 U14380 ( .A0(\xArray[5][37] ), .A1(n8282), .B0(\xArray[9][37] ), 
        .B1(n8228), .C0(n1632), .Y(n1107) );
  OA22X1 U14381 ( .A0(\xArray[1][37] ), .A1(n8200), .B0(\xArray[13][37] ), 
        .B1(n8273), .Y(n1632) );
  OAI221XL U14382 ( .A0(\xArray[9][34] ), .A1(n8291), .B0(\xArray[13][34] ), 
        .B1(n8237), .C0(n873), .Y(n502) );
  OAI221XL U14383 ( .A0(\xArray[9][35] ), .A1(n8291), .B0(\xArray[13][35] ), 
        .B1(n8237), .C0(n870), .Y(n494) );
  OAI221XL U14384 ( .A0(\xArray[2][33] ), .A1(n8288), .B0(\xArray[6][33] ), 
        .B1(n8234), .C0(n2023), .Y(n1643) );
  OAI222XL U14385 ( .A0(n581), .A1(n8339), .B0(n582), .B1(n8309), .C0(n583), 
        .C1(n7730), .Y(n576) );
  AOI221XL U14386 ( .A0(\xArray[14][24] ), .A1(n6573), .B0(\xArray[2][24] ), 
        .B1(n8360), .C0(n578), .Y(n577) );
  OAI22XL U14387 ( .A0(n8359), .A1(n9203), .B0(n6597), .B1(n9205), .Y(n578) );
  MX4X1 U14388 ( .A(n6848), .B(n6846), .C(n6847), .D(n6845), .S0(n7006), .S1(
        n7004), .Y(N25569) );
  MX4X1 U14389 ( .A(n6844), .B(n6842), .C(n6843), .D(n6841), .S0(n7006), .S1(
        n7004), .Y(N25570) );
  MX4X1 U14390 ( .A(\bArray[0][28] ), .B(\bArray[1][28] ), .C(\bArray[2][28] ), 
        .D(\bArray[3][28] ), .S0(n7209), .S1(n7221), .Y(n7059) );
  MX4X1 U14391 ( .A(\bArray[0][31] ), .B(\bArray[1][31] ), .C(\bArray[2][31] ), 
        .D(\bArray[3][31] ), .S0(n7202), .S1(n8409), .Y(n7071) );
  OAI221X1 U14392 ( .A0(\xArray[3][35] ), .A1(n8283), .B0(\xArray[7][35] ), 
        .B1(n8235), .C0(n2007), .Y(n1410) );
  OA22X1 U14393 ( .A0(\xArray[15][35] ), .A1(n8192), .B0(\xArray[11][35] ), 
        .B1(n8265), .Y(n2007) );
  OAI221X1 U14394 ( .A0(\xArray[3][36] ), .A1(n8283), .B0(\xArray[7][36] ), 
        .B1(n8235), .C0(n1998), .Y(n1406) );
  OAI221X1 U14395 ( .A0(\xArray[3][37] ), .A1(n8280), .B0(\xArray[7][37] ), 
        .B1(n8235), .C0(n1989), .Y(n1402) );
  AOI221XL U14396 ( .A0(\xArray[13][28] ), .A1(n8181), .B0(\xArray[1][28] ), 
        .B1(n8178), .C0(n2065), .Y(n2064) );
  OAI22XL U14397 ( .A0(n8174), .A1(n9172), .B0(n8171), .B1(n9170), .Y(n2065)
         );
  AOI221XL U14398 ( .A0(\xArray[13][29] ), .A1(n8179), .B0(\xArray[1][29] ), 
        .B1(n8176), .C0(n2056), .Y(n2055) );
  OAI22XL U14399 ( .A0(n8174), .A1(n9164), .B0(n8171), .B1(n9162), .Y(n2056)
         );
  AOI221XL U14400 ( .A0(\xArray[13][30] ), .A1(n8181), .B0(\xArray[1][30] ), 
        .B1(n8177), .C0(n2047), .Y(n2046) );
  OAI22XL U14401 ( .A0(n8174), .A1(n9156), .B0(n8171), .B1(n9154), .Y(n2047)
         );
  AOI221XL U14402 ( .A0(\xArray[13][31] ), .A1(n8181), .B0(\xArray[1][31] ), 
        .B1(n8177), .C0(n2038), .Y(n2037) );
  OAI22XL U14403 ( .A0(n8174), .A1(n9148), .B0(n8171), .B1(n9146), .Y(n2038)
         );
  OAI221X1 U14404 ( .A0(\xArray[7][37] ), .A1(n8290), .B0(\xArray[11][37] ), 
        .B1(n8226), .C0(n1109), .Y(n477) );
  OAI221X1 U14405 ( .A0(\xArray[7][38] ), .A1(n8284), .B0(\xArray[11][38] ), 
        .B1(n8227), .C0(n1104), .Y(n469) );
  AOI2BB2X1 U14406 ( .B0(n9088), .B1(n8213), .A0N(\xArray[15][38] ), .A1N(
        n8256), .Y(n1104) );
  OAI221X1 U14407 ( .A0(\xArray[4][38] ), .A1(n8283), .B0(\xArray[8][38] ), 
        .B1(n8238), .C0(n1981), .Y(n1396) );
  OAI221X1 U14408 ( .A0(\xArray[4][39] ), .A1(n8280), .B0(\xArray[8][39] ), 
        .B1(n8241), .C0(n1972), .Y(n1392) );
  OAI221X1 U14409 ( .A0(\xArray[8][36] ), .A1(n8292), .B0(\xArray[12][36] ), 
        .B1(n8226), .C0(n1113), .Y(n487) );
  OAI221X1 U14410 ( .A0(\xArray[8][37] ), .A1(n8286), .B0(\xArray[12][37] ), 
        .B1(n8236), .C0(n1108), .Y(n479) );
  OAI221X1 U14411 ( .A0(\xArray[6][37] ), .A1(n8294), .B0(\xArray[10][37] ), 
        .B1(n8240), .C0(n1403), .Y(n863) );
  OAI221X1 U14412 ( .A0(\xArray[6][38] ), .A1(n8294), .B0(\xArray[10][38] ), 
        .B1(n8240), .C0(n1399), .Y(n860) );
  OAI221X1 U14413 ( .A0(\xArray[5][38] ), .A1(n8282), .B0(\xArray[9][38] ), 
        .B1(n8228), .C0(n1629), .Y(n1102) );
  OA22X1 U14414 ( .A0(\xArray[1][38] ), .A1(n8200), .B0(\xArray[13][38] ), 
        .B1(n8273), .Y(n1629) );
  OAI221X1 U14415 ( .A0(\xArray[5][39] ), .A1(n8282), .B0(\xArray[9][39] ), 
        .B1(n8228), .C0(n1626), .Y(n1097) );
  OA22X1 U14416 ( .A0(\xArray[1][39] ), .A1(n8200), .B0(\xArray[13][39] ), 
        .B1(n8270), .Y(n1626) );
  OAI221XL U14417 ( .A0(\xArray[9][36] ), .A1(n8291), .B0(\xArray[13][36] ), 
        .B1(n8237), .C0(n867), .Y(n486) );
  OAI221XL U14418 ( .A0(\xArray[9][37] ), .A1(n8285), .B0(\xArray[13][37] ), 
        .B1(n8232), .C0(n864), .Y(n478) );
  OA22X1 U14419 ( .A0(\xArray[5][37] ), .A1(n8194), .B0(\xArray[1][37] ), .B1(
        n8267), .Y(n864) );
  OAI221XL U14420 ( .A0(\xArray[2][34] ), .A1(n8281), .B0(\xArray[6][34] ), 
        .B1(n8235), .C0(n2014), .Y(n1640) );
  AOI2BB2X1 U14421 ( .B0(n9126), .B1(n8202), .A0N(\xArray[10][34] ), .A1N(
        n8255), .Y(n2014) );
  OAI221XL U14422 ( .A0(\xArray[2][35] ), .A1(n8283), .B0(\xArray[6][35] ), 
        .B1(n8235), .C0(n2005), .Y(n1637) );
  OAI221XL U14423 ( .A0(\xArray[2][36] ), .A1(n8283), .B0(\xArray[6][36] ), 
        .B1(n8235), .C0(n1996), .Y(n1634) );
  OAI222XL U14424 ( .A0(n557), .A1(n8339), .B0(n558), .B1(n8309), .C0(n559), 
        .C1(n7714), .Y(n552) );
  AOI221XL U14425 ( .A0(\xArray[14][27] ), .A1(n6573), .B0(\xArray[2][27] ), 
        .B1(n8360), .C0(n554), .Y(n553) );
  OAI22XL U14426 ( .A0(n8358), .A1(n9179), .B0(n8353), .B1(n9181), .Y(n554) );
  OAI222XL U14427 ( .A0(n565), .A1(n8339), .B0(n566), .B1(n8309), .C0(n567), 
        .C1(n7737), .Y(n560) );
  AOI221XL U14428 ( .A0(\xArray[14][26] ), .A1(n6573), .B0(\xArray[2][26] ), 
        .B1(n8360), .C0(n562), .Y(n561) );
  OAI22XL U14429 ( .A0(n8358), .A1(n9187), .B0(n8353), .B1(n9189), .Y(n562) );
  OAI222XL U14430 ( .A0(n573), .A1(n8339), .B0(n574), .B1(n8309), .C0(n575), 
        .C1(n7717), .Y(n568) );
  AOI221XL U14431 ( .A0(\xArray[14][25] ), .A1(n6573), .B0(\xArray[2][25] ), 
        .B1(n8360), .C0(n570), .Y(n569) );
  OAI22XL U14432 ( .A0(n8358), .A1(n9195), .B0(n8353), .B1(n9197), .Y(n570) );
  MX4X1 U14433 ( .A(n6856), .B(n6854), .C(n6855), .D(n6853), .S0(n7006), .S1(
        n7004), .Y(N25567) );
  MX4X1 U14434 ( .A(n6852), .B(n6850), .C(n6851), .D(n6849), .S0(n7006), .S1(
        n7004), .Y(N25568) );
  OAI221X1 U14435 ( .A0(\xArray[3][38] ), .A1(n8283), .B0(\xArray[7][38] ), 
        .B1(n8238), .C0(n1980), .Y(n1398) );
  OAI221X1 U14436 ( .A0(\xArray[7][39] ), .A1(n8290), .B0(\xArray[11][39] ), 
        .B1(n8227), .C0(n1099), .Y(n461) );
  OAI221X1 U14437 ( .A0(\xArray[4][40] ), .A1(n8280), .B0(\xArray[8][40] ), 
        .B1(n8232), .C0(n1963), .Y(n1388) );
  OAI221X1 U14438 ( .A0(\xArray[4][41] ), .A1(n8295), .B0(\xArray[8][41] ), 
        .B1(n8226), .C0(n1954), .Y(n1384) );
  OAI221X1 U14439 ( .A0(\xArray[8][38] ), .A1(n8284), .B0(\xArray[12][38] ), 
        .B1(n8227), .C0(n1103), .Y(n471) );
  OA22X1 U14440 ( .A0(\xArray[4][38] ), .A1(n8197), .B0(\xArray[0][38] ), .B1(
        n8261), .Y(n1103) );
  OAI221X1 U14441 ( .A0(\xArray[8][39] ), .A1(n8281), .B0(\xArray[12][39] ), 
        .B1(n8227), .C0(n1098), .Y(n463) );
  OAI221X1 U14442 ( .A0(\xArray[6][39] ), .A1(n8294), .B0(\xArray[10][39] ), 
        .B1(n8240), .C0(n1395), .Y(n857) );
  OAI221X1 U14443 ( .A0(\xArray[6][40] ), .A1(n8294), .B0(\xArray[10][40] ), 
        .B1(n8240), .C0(n1391), .Y(n854) );
  OAI221X1 U14444 ( .A0(\xArray[5][40] ), .A1(n8282), .B0(\xArray[9][40] ), 
        .B1(n8228), .C0(n1623), .Y(n1092) );
  OA22X1 U14445 ( .A0(\xArray[1][40] ), .A1(n8199), .B0(\xArray[13][40] ), 
        .B1(n8273), .Y(n1623) );
  OAI221X1 U14446 ( .A0(\xArray[5][41] ), .A1(n8281), .B0(\xArray[9][41] ), 
        .B1(n8225), .C0(n1620), .Y(n1087) );
  OA22X1 U14447 ( .A0(\xArray[1][41] ), .A1(n8199), .B0(\xArray[13][41] ), 
        .B1(n8254), .Y(n1620) );
  OAI221XL U14448 ( .A0(\xArray[9][38] ), .A1(n8296), .B0(\xArray[13][38] ), 
        .B1(n8232), .C0(n861), .Y(n470) );
  OA22X1 U14449 ( .A0(\xArray[5][38] ), .A1(n8194), .B0(\xArray[1][38] ), .B1(
        n8267), .Y(n861) );
  OAI221XL U14450 ( .A0(\xArray[9][39] ), .A1(n8296), .B0(\xArray[13][39] ), 
        .B1(n8232), .C0(n858), .Y(n462) );
  OAI221XL U14451 ( .A0(\xArray[2][37] ), .A1(n8283), .B0(\xArray[6][37] ), 
        .B1(n8235), .C0(n1987), .Y(n1631) );
  OAI221XL U14452 ( .A0(\xArray[2][38] ), .A1(n8280), .B0(\xArray[6][38] ), 
        .B1(n8238), .C0(n1978), .Y(n1628) );
  OAI222XL U14453 ( .A0(n549), .A1(n8339), .B0(n550), .B1(n8309), .C0(n551), 
        .C1(n7737), .Y(n544) );
  AOI221XL U14454 ( .A0(\xArray[14][28] ), .A1(n6573), .B0(\xArray[2][28] ), 
        .B1(n8361), .C0(n546), .Y(n545) );
  OAI22XL U14455 ( .A0(n8358), .A1(n9171), .B0(n8355), .B1(n9173), .Y(n546) );
  MX4X1 U14456 ( .A(n6864), .B(n6862), .C(n6863), .D(n6861), .S0(n7006), .S1(
        n7004), .Y(N25565) );
  MX4X1 U14457 ( .A(n6860), .B(n6858), .C(n6859), .D(n6857), .S0(n7006), .S1(
        n7004), .Y(N25566) );
  OAI221X1 U14458 ( .A0(\xArray[3][39] ), .A1(n8280), .B0(\xArray[7][39] ), 
        .B1(n8238), .C0(n1971), .Y(n1394) );
  OAI221X1 U14459 ( .A0(\xArray[3][40] ), .A1(n8283), .B0(\xArray[7][40] ), 
        .B1(n8238), .C0(n1962), .Y(n1390) );
  AOI221XL U14460 ( .A0(\xArray[13][32] ), .A1(n8181), .B0(\xArray[1][32] ), 
        .B1(n8177), .C0(n2029), .Y(n2028) );
  OAI22XL U14461 ( .A0(n8174), .A1(n9140), .B0(n1751), .B1(n9138), .Y(n2029)
         );
  AOI221XL U14462 ( .A0(\xArray[13][33] ), .A1(n8181), .B0(\xArray[1][33] ), 
        .B1(n8177), .C0(n2020), .Y(n2019) );
  OAI22XL U14463 ( .A0(n8174), .A1(n9132), .B0(n1751), .B1(n9130), .Y(n2020)
         );
  AOI221XL U14464 ( .A0(\xArray[13][34] ), .A1(n8181), .B0(\xArray[1][34] ), 
        .B1(n8177), .C0(n2011), .Y(n2010) );
  OAI22XL U14465 ( .A0(n8173), .A1(n9124), .B0(n1751), .B1(n9122), .Y(n2011)
         );
  AOI221XL U14466 ( .A0(\xArray[13][35] ), .A1(n8180), .B0(\xArray[1][35] ), 
        .B1(n8177), .C0(n2002), .Y(n2001) );
  OAI22XL U14467 ( .A0(n8173), .A1(n9116), .B0(n1751), .B1(n9114), .Y(n2002)
         );
  OAI221X1 U14468 ( .A0(\xArray[7][40] ), .A1(n8281), .B0(\xArray[11][40] ), 
        .B1(n8227), .C0(n1094), .Y(n453) );
  OAI221X1 U14469 ( .A0(\xArray[7][41] ), .A1(n8290), .B0(\xArray[11][41] ), 
        .B1(n8227), .C0(n1089), .Y(n445) );
  OAI221X1 U14470 ( .A0(\xArray[4][42] ), .A1(n8286), .B0(\xArray[8][42] ), 
        .B1(n8236), .C0(n1945), .Y(n1380) );
  OAI221X1 U14471 ( .A0(\xArray[4][43] ), .A1(n8279), .B0(\xArray[8][43] ), 
        .B1(n8225), .C0(n1936), .Y(n1376) );
  OAI221X1 U14472 ( .A0(\xArray[8][40] ), .A1(n8290), .B0(\xArray[12][40] ), 
        .B1(n8227), .C0(n1093), .Y(n455) );
  OAI221X1 U14473 ( .A0(\xArray[8][41] ), .A1(n8290), .B0(\xArray[12][41] ), 
        .B1(n8227), .C0(n1088), .Y(n447) );
  OAI221X1 U14474 ( .A0(\xArray[6][41] ), .A1(n8294), .B0(\xArray[10][41] ), 
        .B1(n8240), .C0(n1387), .Y(n851) );
  OAI221X1 U14475 ( .A0(\xArray[6][42] ), .A1(n8294), .B0(\xArray[10][42] ), 
        .B1(n8240), .C0(n1383), .Y(n848) );
  OAI221X1 U14476 ( .A0(\xArray[5][42] ), .A1(n8281), .B0(\xArray[9][42] ), 
        .B1(n8227), .C0(n1617), .Y(n1082) );
  OAI221XL U14477 ( .A0(\xArray[9][40] ), .A1(n8279), .B0(\xArray[13][40] ), 
        .B1(n8232), .C0(n855), .Y(n454) );
  OAI221XL U14478 ( .A0(\xArray[2][39] ), .A1(n8283), .B0(\xArray[6][39] ), 
        .B1(n8241), .C0(n1969), .Y(n1625) );
  OAI221XL U14479 ( .A0(\xArray[2][40] ), .A1(n8292), .B0(\xArray[6][40] ), 
        .B1(n8236), .C0(n1960), .Y(n1622) );
  OAI222XL U14480 ( .A0(n525), .A1(n8338), .B0(n526), .B1(n8318), .C0(n527), 
        .C1(n7737), .Y(n520) );
  AOI221XL U14481 ( .A0(\xArray[14][31] ), .A1(n6573), .B0(\xArray[2][31] ), 
        .B1(n8360), .C0(n522), .Y(n521) );
  OAI22XL U14482 ( .A0(n8358), .A1(n9147), .B0(n6597), .B1(n9149), .Y(n522) );
  OAI222XL U14483 ( .A0(n533), .A1(n8338), .B0(n534), .B1(n8309), .C0(n535), 
        .C1(n7737), .Y(n528) );
  AOI221XL U14484 ( .A0(\xArray[14][30] ), .A1(n6573), .B0(\xArray[2][30] ), 
        .B1(n8360), .C0(n530), .Y(n529) );
  OAI22XL U14485 ( .A0(n8358), .A1(n9155), .B0(n6597), .B1(n9157), .Y(n530) );
  OAI222XL U14486 ( .A0(n541), .A1(n8339), .B0(n542), .B1(n8309), .C0(n543), 
        .C1(n7737), .Y(n536) );
  AOI221XL U14487 ( .A0(\xArray[14][29] ), .A1(n6573), .B0(\xArray[2][29] ), 
        .B1(n8360), .C0(n538), .Y(n537) );
  OAI22XL U14488 ( .A0(n8358), .A1(n9163), .B0(n6597), .B1(n9165), .Y(n538) );
  MX4X1 U14489 ( .A(n6876), .B(n6874), .C(n6875), .D(n6873), .S0(n7005), .S1(
        n7003), .Y(N25562) );
  MX4X1 U14490 ( .A(n6872), .B(n6870), .C(n6871), .D(n6869), .S0(n7006), .S1(
        n7004), .Y(N25563) );
  MX4X1 U14491 ( .A(n6868), .B(n6866), .C(n6867), .D(n6865), .S0(n7006), .S1(
        n7004), .Y(N25564) );
  OAI221X1 U14492 ( .A0(\xArray[3][41] ), .A1(n8286), .B0(\xArray[7][41] ), 
        .B1(n8226), .C0(n1953), .Y(n1386) );
  OAI221X1 U14493 ( .A0(\xArray[3][42] ), .A1(n8292), .B0(\xArray[7][42] ), 
        .B1(n8226), .C0(n1944), .Y(n1382) );
  AOI221XL U14494 ( .A0(\xArray[13][36] ), .A1(n8180), .B0(\xArray[1][36] ), 
        .B1(n8176), .C0(n1993), .Y(n1992) );
  OAI22XL U14495 ( .A0(n1749), .A1(n9108), .B0(n1751), .B1(n9106), .Y(n1993)
         );
  MX4X1 U14496 ( .A(\bArray[12][38] ), .B(\bArray[13][38] ), .C(
        \bArray[14][38] ), .D(\bArray[15][38] ), .S0(n7207), .S1(n7221), .Y(
        n7096) );
  MX4X1 U14497 ( .A(\bArray[8][38] ), .B(\bArray[9][38] ), .C(\bArray[10][38] ), .D(\bArray[11][38] ), .S0(n7206), .S1(n7221), .Y(n7097) );
  MX4X1 U14498 ( .A(\bArray[4][38] ), .B(\bArray[5][38] ), .C(\bArray[6][38] ), 
        .D(\bArray[7][38] ), .S0(n7206), .S1(n7219), .Y(n7098) );
  OAI221X1 U14499 ( .A0(\xArray[7][42] ), .A1(n8290), .B0(\xArray[11][42] ), 
        .B1(n8235), .C0(n1084), .Y(n437) );
  OAI221X1 U14500 ( .A0(\xArray[7][43] ), .A1(n8290), .B0(\xArray[11][43] ), 
        .B1(n8235), .C0(n1079), .Y(n429) );
  OAI221X1 U14501 ( .A0(\xArray[7][44] ), .A1(n8290), .B0(\xArray[11][44] ), 
        .B1(n8235), .C0(n1074), .Y(n421) );
  OAI221X1 U14502 ( .A0(\xArray[4][44] ), .A1(n8279), .B0(\xArray[8][44] ), 
        .B1(n8225), .C0(n1927), .Y(n1372) );
  OAI221X1 U14503 ( .A0(\xArray[8][42] ), .A1(n8290), .B0(\xArray[12][42] ), 
        .B1(n8235), .C0(n1083), .Y(n439) );
  OAI221X1 U14504 ( .A0(\xArray[8][43] ), .A1(n8290), .B0(\xArray[12][43] ), 
        .B1(n8235), .C0(n1078), .Y(n431) );
  OAI221X1 U14505 ( .A0(\xArray[8][44] ), .A1(n8290), .B0(\xArray[12][44] ), 
        .B1(n8235), .C0(n1073), .Y(n423) );
  OAI221X1 U14506 ( .A0(\xArray[6][43] ), .A1(n8294), .B0(\xArray[10][43] ), 
        .B1(n8240), .C0(n1379), .Y(n845) );
  OAI221X1 U14507 ( .A0(\xArray[6][44] ), .A1(n8294), .B0(\xArray[10][44] ), 
        .B1(n8240), .C0(n1375), .Y(n842) );
  OAI221X1 U14508 ( .A0(\xArray[5][43] ), .A1(n8286), .B0(\xArray[9][43] ), 
        .B1(n8225), .C0(n1614), .Y(n1077) );
  OAI221X1 U14509 ( .A0(\xArray[5][44] ), .A1(n8286), .B0(\xArray[9][44] ), 
        .B1(n8227), .C0(n1611), .Y(n1072) );
  OAI221XL U14510 ( .A0(\xArray[9][41] ), .A1(n8279), .B0(\xArray[13][41] ), 
        .B1(n8232), .C0(n852), .Y(n446) );
  OAI221XL U14511 ( .A0(\xArray[9][42] ), .A1(n8281), .B0(\xArray[13][42] ), 
        .B1(n8232), .C0(n849), .Y(n438) );
  OAI221XL U14512 ( .A0(\xArray[2][41] ), .A1(n8290), .B0(\xArray[6][41] ), 
        .B1(n8236), .C0(n1951), .Y(n1619) );
  OAI221XL U14513 ( .A0(\xArray[2][42] ), .A1(n8279), .B0(\xArray[6][42] ), 
        .B1(n8225), .C0(n1942), .Y(n1616) );
  OAI222XL U14514 ( .A0(n509), .A1(n8338), .B0(n510), .B1(n8309), .C0(n511), 
        .C1(n7737), .Y(n504) );
  AOI221XL U14515 ( .A0(\xArray[14][33] ), .A1(n6573), .B0(\xArray[2][33] ), 
        .B1(n8360), .C0(n506), .Y(n505) );
  OAI22XL U14516 ( .A0(n8358), .A1(n9131), .B0(n6597), .B1(n9133), .Y(n506) );
  OAI222XL U14517 ( .A0(n517), .A1(n8338), .B0(n518), .B1(n8309), .C0(n519), 
        .C1(n7737), .Y(n512) );
  AOI221XL U14518 ( .A0(\xArray[14][32] ), .A1(n6573), .B0(\xArray[2][32] ), 
        .B1(n8360), .C0(n514), .Y(n513) );
  OAI22XL U14519 ( .A0(n8358), .A1(n9139), .B0(n6597), .B1(n9141), .Y(n514) );
  MX4X1 U14520 ( .A(n6880), .B(n6878), .C(n6879), .D(n6877), .S0(n8411), .S1(
        n7004), .Y(N25561) );
  MX4X1 U14521 ( .A(\bArray[8][39] ), .B(\bArray[9][39] ), .C(\bArray[10][39] ), .D(\bArray[11][39] ), .S0(n6984), .S1(n6994), .Y(n6878) );
  MX4X1 U14522 ( .A(\bArray[0][39] ), .B(\bArray[1][39] ), .C(\bArray[2][39] ), 
        .D(\bArray[3][39] ), .S0(n6980), .S1(n6995), .Y(n6880) );
  MX4X1 U14523 ( .A(\bArray[12][39] ), .B(\bArray[13][39] ), .C(
        \bArray[14][39] ), .D(\bArray[15][39] ), .S0(n6979), .S1(n6994), .Y(
        n6877) );
  MX4X1 U14524 ( .A(\bArray[4][39] ), .B(\bArray[5][39] ), .C(\bArray[6][39] ), 
        .D(\bArray[7][39] ), .S0(n6979), .S1(n6995), .Y(n6879) );
  MX4X1 U14525 ( .A(\bArray[0][38] ), .B(\bArray[1][38] ), .C(\bArray[2][38] ), 
        .D(\bArray[3][38] ), .S0(n7207), .S1(n7221), .Y(n7099) );
  OAI221X1 U14526 ( .A0(\xArray[3][43] ), .A1(n8279), .B0(\xArray[7][43] ), 
        .B1(n8225), .C0(n1935), .Y(n1378) );
  AOI221XL U14527 ( .A0(\xArray[13][37] ), .A1(n8180), .B0(\xArray[1][37] ), 
        .B1(n8176), .C0(n1984), .Y(n1983) );
  OAI22XL U14528 ( .A0(n8173), .A1(n9100), .B0(n8171), .B1(n9098), .Y(n1984)
         );
  AOI221XL U14529 ( .A0(\xArray[13][38] ), .A1(n8180), .B0(\xArray[1][38] ), 
        .B1(n8176), .C0(n1975), .Y(n1974) );
  OAI22XL U14530 ( .A0(n8174), .A1(n9092), .B0(n8171), .B1(n9090), .Y(n1975)
         );
  AOI221XL U14531 ( .A0(\xArray[13][39] ), .A1(n8180), .B0(\xArray[1][39] ), 
        .B1(n8176), .C0(n1966), .Y(n1965) );
  OAI22XL U14532 ( .A0(n8174), .A1(n9084), .B0(n8170), .B1(n9082), .Y(n1966)
         );
  OAI221X1 U14533 ( .A0(\xArray[7][45] ), .A1(n8290), .B0(\xArray[11][45] ), 
        .B1(n8235), .C0(n1069), .Y(n413) );
  OAI221X1 U14534 ( .A0(\xArray[7][46] ), .A1(n8290), .B0(\xArray[11][46] ), 
        .B1(n8235), .C0(n1064), .Y(n405) );
  OAI221X1 U14535 ( .A0(\xArray[4][45] ), .A1(n8279), .B0(\xArray[8][45] ), 
        .B1(n8225), .C0(n1918), .Y(n1368) );
  OAI221X1 U14536 ( .A0(\xArray[4][46] ), .A1(n8279), .B0(\xArray[8][46] ), 
        .B1(n8225), .C0(n1909), .Y(n1364) );
  OAI221X1 U14537 ( .A0(\xArray[4][47] ), .A1(n8279), .B0(\xArray[8][47] ), 
        .B1(n8225), .C0(n1900), .Y(n1360) );
  OAI221X1 U14538 ( .A0(\xArray[8][45] ), .A1(n8290), .B0(\xArray[12][45] ), 
        .B1(n8235), .C0(n1068), .Y(n415) );
  OAI221X1 U14539 ( .A0(\xArray[6][45] ), .A1(n8294), .B0(\xArray[10][45] ), 
        .B1(n8240), .C0(n1371), .Y(n839) );
  OAI221X1 U14540 ( .A0(\xArray[6][46] ), .A1(n8279), .B0(\xArray[10][46] ), 
        .B1(n8233), .C0(n1367), .Y(n836) );
  OAI221X1 U14541 ( .A0(\xArray[5][45] ), .A1(n8281), .B0(\xArray[9][45] ), 
        .B1(n8227), .C0(n1608), .Y(n1067) );
  OAI221X1 U14542 ( .A0(\xArray[5][46] ), .A1(n8286), .B0(\xArray[9][46] ), 
        .B1(n8227), .C0(n1605), .Y(n1062) );
  OAI221X1 U14543 ( .A0(\xArray[5][47] ), .A1(n8286), .B0(\xArray[9][47] ), 
        .B1(n8225), .C0(n1602), .Y(n1057) );
  OAI221XL U14544 ( .A0(\xArray[9][43] ), .A1(n8281), .B0(\xArray[13][43] ), 
        .B1(n8232), .C0(n846), .Y(n430) );
  OAI221XL U14545 ( .A0(\xArray[9][44] ), .A1(n8281), .B0(\xArray[13][44] ), 
        .B1(n8232), .C0(n843), .Y(n422) );
  OAI221XL U14546 ( .A0(\xArray[2][43] ), .A1(n8279), .B0(\xArray[6][43] ), 
        .B1(n8225), .C0(n1933), .Y(n1613) );
  OAI222XL U14547 ( .A0(n493), .A1(n8338), .B0(n494), .B1(n8318), .C0(n495), 
        .C1(n7713), .Y(n488) );
  AOI221XL U14548 ( .A0(\xArray[14][35] ), .A1(n6573), .B0(\xArray[2][35] ), 
        .B1(n8360), .C0(n490), .Y(n489) );
  OAI22XL U14549 ( .A0(n8358), .A1(n9115), .B0(n8353), .B1(n9117), .Y(n490) );
  OAI222XL U14550 ( .A0(n501), .A1(n8338), .B0(n502), .B1(n8309), .C0(n503), 
        .C1(n7737), .Y(n496) );
  AOI221XL U14551 ( .A0(\xArray[14][34] ), .A1(n6573), .B0(\xArray[2][34] ), 
        .B1(n8360), .C0(n498), .Y(n497) );
  OAI22XL U14552 ( .A0(n8358), .A1(n9123), .B0(n8353), .B1(n9125), .Y(n498) );
  MX4X1 U14553 ( .A(n6892), .B(n6890), .C(n6891), .D(n6889), .S0(N1760), .S1(
        n8412), .Y(N25558) );
  MX4X1 U14554 ( .A(\bArray[8][42] ), .B(\bArray[9][42] ), .C(\bArray[10][42] ), .D(\bArray[11][42] ), .S0(n6980), .S1(n6992), .Y(n6890) );
  MX4X1 U14555 ( .A(\bArray[0][42] ), .B(\bArray[1][42] ), .C(\bArray[2][42] ), 
        .D(\bArray[3][42] ), .S0(n6980), .S1(n6992), .Y(n6892) );
  MX4X1 U14556 ( .A(\bArray[12][42] ), .B(\bArray[13][42] ), .C(
        \bArray[14][42] ), .D(\bArray[15][42] ), .S0(n6980), .S1(n6992), .Y(
        n6889) );
  MX4X1 U14557 ( .A(n6888), .B(n6886), .C(n6887), .D(n6885), .S0(N1760), .S1(
        N1759), .Y(N25559) );
  MX4X1 U14558 ( .A(\bArray[8][41] ), .B(\bArray[9][41] ), .C(\bArray[10][41] ), .D(\bArray[11][41] ), .S0(n6979), .S1(n6992), .Y(n6886) );
  MX4X1 U14559 ( .A(\bArray[0][41] ), .B(\bArray[1][41] ), .C(\bArray[2][41] ), 
        .D(\bArray[3][41] ), .S0(n6984), .S1(n6998), .Y(n6888) );
  MX4X1 U14560 ( .A(\bArray[12][41] ), .B(\bArray[13][41] ), .C(
        \bArray[14][41] ), .D(\bArray[15][41] ), .S0(n6979), .S1(n8413), .Y(
        n6885) );
  MX4X1 U14561 ( .A(n6884), .B(n6882), .C(n6883), .D(n6881), .S0(N1760), .S1(
        n8412), .Y(N25560) );
  MX4X1 U14562 ( .A(\bArray[8][40] ), .B(\bArray[9][40] ), .C(\bArray[10][40] ), .D(\bArray[11][40] ), .S0(n6979), .S1(n8413), .Y(n6882) );
  MX4X1 U14563 ( .A(\bArray[0][40] ), .B(\bArray[1][40] ), .C(\bArray[2][40] ), 
        .D(\bArray[3][40] ), .S0(n6980), .S1(n6995), .Y(n6884) );
  MX4X1 U14564 ( .A(\bArray[12][40] ), .B(\bArray[13][40] ), .C(
        \bArray[14][40] ), .D(\bArray[15][40] ), .S0(n6979), .S1(n6995), .Y(
        n6881) );
  CLKINVX1 U14565 ( .A(\xArray[14][42] ), .Y(n9062) );
  CLKINVX1 U14566 ( .A(\xArray[3][42] ), .Y(n9056) );
  CLKINVX1 U14567 ( .A(\xArray[3][43] ), .Y(n9048) );
  CLKINVX1 U14568 ( .A(\xArray[3][44] ), .Y(n9040) );
  MX4X1 U14569 ( .A(\bArray[4][42] ), .B(\bArray[5][42] ), .C(\bArray[6][42] ), 
        .D(\bArray[7][42] ), .S0(n6980), .S1(n6991), .Y(n6891) );
  MX4X1 U14570 ( .A(\bArray[4][41] ), .B(\bArray[5][41] ), .C(\bArray[6][41] ), 
        .D(\bArray[7][41] ), .S0(n6979), .S1(n8413), .Y(n6887) );
  MX4X1 U14571 ( .A(\bArray[4][40] ), .B(\bArray[5][40] ), .C(\bArray[6][40] ), 
        .D(\bArray[7][40] ), .S0(n6980), .S1(n6995), .Y(n6883) );
  OAI221X1 U14572 ( .A0(\xArray[3][44] ), .A1(n8279), .B0(\xArray[7][44] ), 
        .B1(n8225), .C0(n1926), .Y(n1374) );
  OAI221X1 U14573 ( .A0(\xArray[3][45] ), .A1(n8279), .B0(\xArray[7][45] ), 
        .B1(n8225), .C0(n1917), .Y(n1370) );
  OAI221X1 U14574 ( .A0(\xArray[3][46] ), .A1(n8279), .B0(\xArray[7][46] ), 
        .B1(n8225), .C0(n1908), .Y(n1366) );
  OAI221X1 U14575 ( .A0(\xArray[3][47] ), .A1(n8279), .B0(\xArray[7][47] ), 
        .B1(n8225), .C0(n1899), .Y(n1362) );
  AOI221XL U14576 ( .A0(\xArray[13][40] ), .A1(n8180), .B0(\xArray[1][40] ), 
        .B1(n8176), .C0(n1957), .Y(n1956) );
  OAI22XL U14577 ( .A0(n8174), .A1(n9076), .B0(n8170), .B1(n9074), .Y(n1957)
         );
  MX4X1 U14578 ( .A(\bArray[8][41] ), .B(\bArray[9][41] ), .C(\bArray[10][41] ), .D(\bArray[11][41] ), .S0(n8410), .S1(n7215), .Y(n7109) );
  MX4X1 U14579 ( .A(\bArray[4][41] ), .B(\bArray[5][41] ), .C(\bArray[6][41] ), 
        .D(\bArray[7][41] ), .S0(n8410), .S1(n7215), .Y(n7110) );
  OAI221X1 U14580 ( .A0(\xArray[7][47] ), .A1(n8287), .B0(\xArray[11][47] ), 
        .B1(n8242), .C0(n1059), .Y(n397) );
  OAI221X1 U14581 ( .A0(\xArray[7][48] ), .A1(n8287), .B0(\xArray[11][48] ), 
        .B1(n8242), .C0(n1054), .Y(n389) );
  OAI221X1 U14582 ( .A0(\xArray[4][48] ), .A1(n8279), .B0(\xArray[8][48] ), 
        .B1(n8234), .C0(n1891), .Y(n1356) );
  OAI221X1 U14583 ( .A0(\xArray[4][49] ), .A1(n8281), .B0(\xArray[8][49] ), 
        .B1(n8226), .C0(n1882), .Y(n1352) );
  OAI221X1 U14584 ( .A0(\xArray[8][46] ), .A1(n8290), .B0(\xArray[12][46] ), 
        .B1(n8235), .C0(n1063), .Y(n407) );
  OAI221X1 U14585 ( .A0(\xArray[8][47] ), .A1(n8287), .B0(\xArray[12][47] ), 
        .B1(n8242), .C0(n1058), .Y(n399) );
  OAI221X1 U14586 ( .A0(\xArray[6][47] ), .A1(n8279), .B0(\xArray[10][47] ), 
        .B1(n8233), .C0(n1363), .Y(n833) );
  OAI221X1 U14587 ( .A0(\xArray[6][48] ), .A1(n8279), .B0(\xArray[10][48] ), 
        .B1(n8233), .C0(n1359), .Y(n830) );
  OAI221X1 U14588 ( .A0(\xArray[5][48] ), .A1(n8292), .B0(\xArray[9][48] ), 
        .B1(n8227), .C0(n1599), .Y(n1052) );
  OAI221X1 U14589 ( .A0(\xArray[5][49] ), .A1(n8286), .B0(\xArray[9][49] ), 
        .B1(n8227), .C0(n1596), .Y(n1047) );
  OAI221XL U14590 ( .A0(\xArray[9][45] ), .A1(n8281), .B0(\xArray[13][45] ), 
        .B1(n8232), .C0(n840), .Y(n414) );
  OAI221XL U14591 ( .A0(\xArray[9][46] ), .A1(n8281), .B0(\xArray[13][46] ), 
        .B1(n8232), .C0(n837), .Y(n406) );
  OAI221XL U14592 ( .A0(\xArray[2][44] ), .A1(n8279), .B0(\xArray[6][44] ), 
        .B1(n8225), .C0(n1924), .Y(n1610) );
  OAI221XL U14593 ( .A0(\xArray[2][45] ), .A1(n8279), .B0(\xArray[6][45] ), 
        .B1(n8225), .C0(n1915), .Y(n1607) );
  OAI221XL U14594 ( .A0(\xArray[2][46] ), .A1(n8279), .B0(\xArray[6][46] ), 
        .B1(n8225), .C0(n1906), .Y(n1604) );
  OAI222XL U14595 ( .A0(n477), .A1(n8338), .B0(n478), .B1(n8314), .C0(n479), 
        .C1(n7733), .Y(n472) );
  AOI221XL U14596 ( .A0(\xArray[14][37] ), .A1(n6573), .B0(\xArray[2][37] ), 
        .B1(n8360), .C0(n474), .Y(n473) );
  OAI22XL U14597 ( .A0(n8358), .A1(n9099), .B0(n8353), .B1(n9101), .Y(n474) );
  OAI222XL U14598 ( .A0(n485), .A1(n8338), .B0(n486), .B1(n8320), .C0(n487), 
        .C1(n7740), .Y(n480) );
  AOI221XL U14599 ( .A0(\xArray[14][36] ), .A1(n6573), .B0(\xArray[2][36] ), 
        .B1(n8360), .C0(n482), .Y(n481) );
  OAI22XL U14600 ( .A0(n8358), .A1(n9107), .B0(n8353), .B1(n9109), .Y(n482) );
  MX4X1 U14601 ( .A(n6896), .B(n6894), .C(n6895), .D(n6893), .S0(n8411), .S1(
        n8412), .Y(N25557) );
  MX4X1 U14602 ( .A(\bArray[8][43] ), .B(\bArray[9][43] ), .C(\bArray[10][43] ), .D(\bArray[11][43] ), .S0(n6980), .S1(n6992), .Y(n6894) );
  MX4X1 U14603 ( .A(\bArray[0][43] ), .B(\bArray[1][43] ), .C(\bArray[2][43] ), 
        .D(\bArray[3][43] ), .S0(n6980), .S1(n6992), .Y(n6896) );
  MX4X1 U14604 ( .A(\bArray[12][43] ), .B(\bArray[13][43] ), .C(
        \bArray[14][43] ), .D(\bArray[15][43] ), .S0(n6980), .S1(n6992), .Y(
        n6893) );
  CLKINVX1 U14605 ( .A(\xArray[14][43] ), .Y(n9054) );
  CLKINVX1 U14606 ( .A(\xArray[14][44] ), .Y(n9046) );
  CLKINVX1 U14607 ( .A(\xArray[3][45] ), .Y(n9032) );
  CLKINVX1 U14608 ( .A(\xArray[3][46] ), .Y(n9024) );
  MX4X1 U14609 ( .A(\bArray[4][43] ), .B(\bArray[5][43] ), .C(\bArray[6][43] ), 
        .D(\bArray[7][43] ), .S0(n6980), .S1(n6992), .Y(n6895) );
  MX4X1 U14610 ( .A(\bArray[0][41] ), .B(\bArray[1][41] ), .C(\bArray[2][41] ), 
        .D(\bArray[3][41] ), .S0(n8410), .S1(n7215), .Y(n7111) );
  OAI221X1 U14611 ( .A0(\xArray[3][48] ), .A1(n8287), .B0(\xArray[7][48] ), 
        .B1(n8240), .C0(n1890), .Y(n1358) );
  OAI221X1 U14612 ( .A0(\xArray[3][49] ), .A1(n8286), .B0(\xArray[7][49] ), 
        .B1(n8224), .C0(n1881), .Y(n1354) );
  AOI221XL U14613 ( .A0(\xArray[13][41] ), .A1(n8181), .B0(\xArray[1][41] ), 
        .B1(n8176), .C0(n1948), .Y(n1947) );
  OAI22XL U14614 ( .A0(n8174), .A1(n9068), .B0(n8170), .B1(n9066), .Y(n1948)
         );
  AOI221XL U14615 ( .A0(\xArray[13][42] ), .A1(n8179), .B0(\xArray[1][42] ), 
        .B1(n8177), .C0(n1939), .Y(n1938) );
  OAI22XL U14616 ( .A0(n8174), .A1(n9060), .B0(n8170), .B1(n9058), .Y(n1939)
         );
  AOI221XL U14617 ( .A0(\xArray[13][43] ), .A1(n8179), .B0(\xArray[1][43] ), 
        .B1(n8177), .C0(n1930), .Y(n1929) );
  OAI22XL U14618 ( .A0(n8174), .A1(n9052), .B0(n8170), .B1(n9050), .Y(n1930)
         );
  MX4X1 U14619 ( .A(\bArray[4][44] ), .B(\bArray[5][44] ), .C(\bArray[6][44] ), 
        .D(\bArray[7][44] ), .S0(n7207), .S1(n7214), .Y(n7122) );
  OAI221X1 U14620 ( .A0(\xArray[7][49] ), .A1(n8287), .B0(\xArray[11][49] ), 
        .B1(n8225), .C0(n1049), .Y(n381) );
  OAI221X1 U14621 ( .A0(\xArray[7][50] ), .A1(n8291), .B0(\xArray[11][50] ), 
        .B1(n8225), .C0(n1044), .Y(n373) );
  OAI221X1 U14622 ( .A0(\xArray[4][50] ), .A1(n8283), .B0(\xArray[8][50] ), 
        .B1(n8233), .C0(n1873), .Y(n1348) );
  OAI221X1 U14623 ( .A0(\xArray[4][51] ), .A1(n8286), .B0(\xArray[8][51] ), 
        .B1(n8233), .C0(n1864), .Y(n1344) );
  OAI221X1 U14624 ( .A0(\xArray[8][48] ), .A1(n8287), .B0(\xArray[12][48] ), 
        .B1(n8242), .C0(n1053), .Y(n391) );
  OAI221X1 U14625 ( .A0(\xArray[8][49] ), .A1(n8287), .B0(\xArray[12][49] ), 
        .B1(n8225), .C0(n1048), .Y(n383) );
  OAI221X1 U14626 ( .A0(\xArray[6][49] ), .A1(n8279), .B0(\xArray[10][49] ), 
        .B1(n8233), .C0(n1355), .Y(n827) );
  OAI221X1 U14627 ( .A0(\xArray[6][50] ), .A1(n8279), .B0(\xArray[10][50] ), 
        .B1(n8233), .C0(n1351), .Y(n824) );
  OAI221X1 U14628 ( .A0(\xArray[5][50] ), .A1(n8292), .B0(\xArray[9][50] ), 
        .B1(n8227), .C0(n1593), .Y(n1042) );
  OAI221X1 U14629 ( .A0(\xArray[5][51] ), .A1(n8295), .B0(\xArray[9][51] ), 
        .B1(n8225), .C0(n1590), .Y(n1037) );
  OAI221XL U14630 ( .A0(\xArray[9][47] ), .A1(n8281), .B0(\xArray[13][47] ), 
        .B1(n8232), .C0(n834), .Y(n398) );
  OAI221XL U14631 ( .A0(\xArray[9][48] ), .A1(n8281), .B0(\xArray[13][48] ), 
        .B1(n8232), .C0(n831), .Y(n390) );
  OAI221XL U14632 ( .A0(\xArray[2][47] ), .A1(n8288), .B0(\xArray[6][47] ), 
        .B1(n8226), .C0(n1897), .Y(n1601) );
  OAI221XL U14633 ( .A0(\xArray[2][48] ), .A1(n8288), .B0(\xArray[6][48] ), 
        .B1(n8234), .C0(n1888), .Y(n1598) );
  OAI222XL U14634 ( .A0(n461), .A1(n8338), .B0(n462), .B1(n8310), .C0(n463), 
        .C1(n7733), .Y(n456) );
  AOI221XL U14635 ( .A0(\xArray[14][39] ), .A1(n6573), .B0(\xArray[2][39] ), 
        .B1(n8362), .C0(n458), .Y(n457) );
  OAI22XL U14636 ( .A0(n8359), .A1(n9083), .B0(n6597), .B1(n9085), .Y(n458) );
  OAI222XL U14637 ( .A0(n469), .A1(n8338), .B0(n470), .B1(n8314), .C0(n471), 
        .C1(n7733), .Y(n464) );
  AOI221XL U14638 ( .A0(\xArray[14][38] ), .A1(n6573), .B0(\xArray[2][38] ), 
        .B1(n8360), .C0(n466), .Y(n465) );
  OAI22XL U14639 ( .A0(n8358), .A1(n9091), .B0(n6597), .B1(n9093), .Y(n466) );
  MX4X1 U14640 ( .A(n6912), .B(n6910), .C(n6911), .D(n6909), .S0(n8411), .S1(
        n8412), .Y(N25553) );
  MX4X1 U14641 ( .A(\bArray[8][47] ), .B(\bArray[9][47] ), .C(\bArray[10][47] ), .D(\bArray[11][47] ), .S0(n6980), .S1(n7001), .Y(n6910) );
  MX4X1 U14642 ( .A(\bArray[0][47] ), .B(\bArray[1][47] ), .C(\bArray[2][47] ), 
        .D(\bArray[3][47] ), .S0(n6983), .S1(n7001), .Y(n6912) );
  MX4X1 U14643 ( .A(\bArray[12][47] ), .B(\bArray[13][47] ), .C(
        \bArray[14][47] ), .D(\bArray[15][47] ), .S0(n6990), .S1(n7001), .Y(
        n6909) );
  MX4X1 U14644 ( .A(n6908), .B(n6906), .C(n6907), .D(n6905), .S0(n8411), .S1(
        n8412), .Y(N25554) );
  MX4X1 U14645 ( .A(\bArray[8][46] ), .B(\bArray[9][46] ), .C(\bArray[10][46] ), .D(\bArray[11][46] ), .S0(n6990), .S1(n7002), .Y(n6906) );
  MX4X1 U14646 ( .A(\bArray[0][46] ), .B(\bArray[1][46] ), .C(\bArray[2][46] ), 
        .D(\bArray[3][46] ), .S0(n6990), .S1(n6992), .Y(n6908) );
  MX4X1 U14647 ( .A(\bArray[12][46] ), .B(\bArray[13][46] ), .C(
        \bArray[14][46] ), .D(\bArray[15][46] ), .S0(n6978), .S1(n7002), .Y(
        n6905) );
  MX4X1 U14648 ( .A(n6904), .B(n6902), .C(n6903), .D(n6901), .S0(n8411), .S1(
        n8412), .Y(N25555) );
  MX4X1 U14649 ( .A(\bArray[8][45] ), .B(\bArray[9][45] ), .C(\bArray[10][45] ), .D(\bArray[11][45] ), .S0(n6987), .S1(n7002), .Y(n6902) );
  MX4X1 U14650 ( .A(\bArray[0][45] ), .B(\bArray[1][45] ), .C(\bArray[2][45] ), 
        .D(\bArray[3][45] ), .S0(n6986), .S1(n7002), .Y(n6904) );
  MX4X1 U14651 ( .A(\bArray[12][45] ), .B(\bArray[13][45] ), .C(
        \bArray[14][45] ), .D(\bArray[15][45] ), .S0(n6988), .S1(n7002), .Y(
        n6901) );
  MX4X1 U14652 ( .A(n6900), .B(n6898), .C(n6899), .D(n6897), .S0(n8411), .S1(
        n8412), .Y(N25556) );
  MX4X1 U14653 ( .A(\bArray[8][44] ), .B(\bArray[9][44] ), .C(\bArray[10][44] ), .D(\bArray[11][44] ), .S0(n6984), .S1(n6992), .Y(n6898) );
  MX4X1 U14654 ( .A(\bArray[0][44] ), .B(\bArray[1][44] ), .C(\bArray[2][44] ), 
        .D(\bArray[3][44] ), .S0(n6987), .S1(n7002), .Y(n6900) );
  MX4X1 U14655 ( .A(\bArray[12][44] ), .B(\bArray[13][44] ), .C(
        \bArray[14][44] ), .D(\bArray[15][44] ), .S0(n6983), .S1(n6992), .Y(
        n6897) );
  CLKINVX1 U14656 ( .A(\xArray[14][45] ), .Y(n9038) );
  CLKINVX1 U14657 ( .A(\xArray[14][46] ), .Y(n9030) );
  CLKINVX1 U14658 ( .A(\xArray[3][47] ), .Y(n9016) );
  CLKINVX1 U14659 ( .A(\xArray[3][48] ), .Y(n9008) );
  MX4X1 U14660 ( .A(\bArray[4][47] ), .B(\bArray[5][47] ), .C(\bArray[6][47] ), 
        .D(\bArray[7][47] ), .S0(n6990), .S1(n6992), .Y(n6911) );
  MX4X1 U14661 ( .A(\bArray[4][46] ), .B(\bArray[5][46] ), .C(\bArray[6][46] ), 
        .D(\bArray[7][46] ), .S0(n6990), .S1(n7002), .Y(n6907) );
  MX4X1 U14662 ( .A(\bArray[4][45] ), .B(\bArray[5][45] ), .C(\bArray[6][45] ), 
        .D(\bArray[7][45] ), .S0(n6987), .S1(n7002), .Y(n6903) );
  MX4X1 U14663 ( .A(\bArray[4][44] ), .B(\bArray[5][44] ), .C(\bArray[6][44] ), 
        .D(\bArray[7][44] ), .S0(n6988), .S1(n8413), .Y(n6899) );
  MX4X1 U14664 ( .A(\bArray[0][44] ), .B(\bArray[1][44] ), .C(\bArray[2][44] ), 
        .D(\bArray[3][44] ), .S0(n7201), .S1(n7222), .Y(n7123) );
  OAI221X1 U14665 ( .A0(\xArray[3][50] ), .A1(n8290), .B0(\xArray[7][50] ), 
        .B1(n8233), .C0(n1872), .Y(n1350) );
  AOI221XL U14666 ( .A0(\xArray[13][44] ), .A1(n8179), .B0(\xArray[1][44] ), 
        .B1(n8177), .C0(n1921), .Y(n1920) );
  OAI22XL U14667 ( .A0(n8174), .A1(n9044), .B0(n8170), .B1(n9042), .Y(n1921)
         );
  MX4X1 U14668 ( .A(\bArray[12][45] ), .B(\bArray[13][45] ), .C(
        \bArray[14][45] ), .D(\bArray[15][45] ), .S0(n7203), .S1(n7213), .Y(
        n7124) );
  MX4X1 U14669 ( .A(\bArray[8][45] ), .B(\bArray[9][45] ), .C(\bArray[10][45] ), .D(\bArray[11][45] ), .S0(n7203), .S1(n7214), .Y(n7125) );
  MX4X1 U14670 ( .A(\bArray[4][45] ), .B(\bArray[5][45] ), .C(\bArray[6][45] ), 
        .D(\bArray[7][45] ), .S0(n7203), .S1(n7214), .Y(n7126) );
  MX4X1 U14671 ( .A(\bArray[12][46] ), .B(\bArray[13][46] ), .C(
        \bArray[14][46] ), .D(\bArray[15][46] ), .S0(n7203), .S1(n7214), .Y(
        n7128) );
  MX4X1 U14672 ( .A(\bArray[8][46] ), .B(\bArray[9][46] ), .C(\bArray[10][46] ), .D(\bArray[11][46] ), .S0(n7203), .S1(n7214), .Y(n7129) );
  MX4X1 U14673 ( .A(\bArray[4][46] ), .B(\bArray[5][46] ), .C(\bArray[6][46] ), 
        .D(\bArray[7][46] ), .S0(n7203), .S1(n7214), .Y(n7130) );
  MX4X1 U14674 ( .A(\bArray[12][47] ), .B(\bArray[13][47] ), .C(
        \bArray[14][47] ), .D(\bArray[15][47] ), .S0(n7203), .S1(n7214), .Y(
        n7132) );
  MX4X1 U14675 ( .A(\bArray[8][47] ), .B(\bArray[9][47] ), .C(\bArray[10][47] ), .D(\bArray[11][47] ), .S0(n7207), .S1(n7221), .Y(n7133) );
  MX4X1 U14676 ( .A(\bArray[4][47] ), .B(\bArray[5][47] ), .C(\bArray[6][47] ), 
        .D(\bArray[7][47] ), .S0(n7207), .S1(N1762), .Y(n7134) );
  OAI221X1 U14677 ( .A0(\xArray[7][51] ), .A1(n8291), .B0(\xArray[11][51] ), 
        .B1(n8225), .C0(n1039), .Y(n365) );
  OAI221X1 U14678 ( .A0(\xArray[4][52] ), .A1(n8286), .B0(\xArray[8][52] ), 
        .B1(n8233), .C0(n1855), .Y(n1340) );
  OAI221X1 U14679 ( .A0(\xArray[8][50] ), .A1(n8282), .B0(\xArray[12][50] ), 
        .B1(n8225), .C0(n1043), .Y(n375) );
  OAI221X1 U14680 ( .A0(\xArray[8][51] ), .A1(n8291), .B0(\xArray[12][51] ), 
        .B1(n8242), .C0(n1038), .Y(n367) );
  OAI221X1 U14681 ( .A0(\xArray[6][51] ), .A1(n8279), .B0(\xArray[10][51] ), 
        .B1(n8228), .C0(n1347), .Y(n821) );
  OAI221X1 U14682 ( .A0(\xArray[6][52] ), .A1(n8279), .B0(\xArray[10][52] ), 
        .B1(n8233), .C0(n1343), .Y(n818) );
  OAI221X1 U14683 ( .A0(\xArray[5][52] ), .A1(n8281), .B0(\xArray[9][52] ), 
        .B1(n8227), .C0(n1587), .Y(n1032) );
  OAI221XL U14684 ( .A0(\xArray[9][49] ), .A1(n8281), .B0(\xArray[13][49] ), 
        .B1(n8238), .C0(n828), .Y(n382) );
  OAI221XL U14685 ( .A0(\xArray[9][50] ), .A1(n8281), .B0(\xArray[13][50] ), 
        .B1(n8232), .C0(n825), .Y(n374) );
  OAI221XL U14686 ( .A0(\xArray[2][49] ), .A1(n8281), .B0(\xArray[6][49] ), 
        .B1(n8226), .C0(n1879), .Y(n1595) );
  OAI221XL U14687 ( .A0(\xArray[2][50] ), .A1(n8281), .B0(\xArray[6][50] ), 
        .B1(n8233), .C0(n1870), .Y(n1592) );
  OAI222XL U14688 ( .A0(n445), .A1(n8338), .B0(n446), .B1(n8310), .C0(n447), 
        .C1(n7707), .Y(n440) );
  AOI221XL U14689 ( .A0(\xArray[14][41] ), .A1(n6573), .B0(\xArray[2][41] ), 
        .B1(n6579), .C0(n442), .Y(n441) );
  OAI22XL U14690 ( .A0(n8356), .A1(n9067), .B0(n8354), .B1(n9069), .Y(n442) );
  OAI222XL U14691 ( .A0(n453), .A1(n8338), .B0(n454), .B1(n8310), .C0(n455), 
        .C1(n7733), .Y(n448) );
  AOI221XL U14692 ( .A0(\xArray[14][40] ), .A1(n6573), .B0(\xArray[2][40] ), 
        .B1(n8362), .C0(n450), .Y(n449) );
  OAI22XL U14693 ( .A0(n8356), .A1(n9075), .B0(n6597), .B1(n9077), .Y(n450) );
  CLKINVX1 U14694 ( .A(\xArray[14][47] ), .Y(n9022) );
  CLKINVX1 U14695 ( .A(\xArray[14][48] ), .Y(n9014) );
  CLKINVX1 U14696 ( .A(\xArray[5][42] ), .Y(n9058) );
  CLKINVX1 U14697 ( .A(\xArray[5][43] ), .Y(n9050) );
  CLKINVX1 U14698 ( .A(\xArray[3][49] ), .Y(n9000) );
  CLKINVX1 U14699 ( .A(\xArray[3][50] ), .Y(n8992) );
  MX4X1 U14700 ( .A(\bArray[0][45] ), .B(\bArray[1][45] ), .C(\bArray[2][45] ), 
        .D(\bArray[3][45] ), .S0(n7207), .S1(n7221), .Y(n7127) );
  MX4X1 U14701 ( .A(\bArray[0][46] ), .B(\bArray[1][46] ), .C(\bArray[2][46] ), 
        .D(\bArray[3][46] ), .S0(n7203), .S1(n7214), .Y(n7131) );
  MX4X1 U14702 ( .A(\bArray[0][47] ), .B(\bArray[1][47] ), .C(\bArray[2][47] ), 
        .D(\bArray[3][47] ), .S0(n7207), .S1(n7214), .Y(n7135) );
  CLKINVX1 U14703 ( .A(\xArray[9][42] ), .Y(n9060) );
  CLKINVX1 U14704 ( .A(\xArray[9][43] ), .Y(n9052) );
  OAI221X1 U14705 ( .A0(\xArray[3][51] ), .A1(n8278), .B0(\xArray[7][51] ), 
        .B1(n8233), .C0(n1863), .Y(n1346) );
  OAI221X1 U14706 ( .A0(\xArray[3][52] ), .A1(n8278), .B0(\xArray[7][52] ), 
        .B1(n8233), .C0(n1854), .Y(n1342) );
  AOI221XL U14707 ( .A0(\xArray[13][45] ), .A1(n8179), .B0(\xArray[1][45] ), 
        .B1(n8177), .C0(n1912), .Y(n1911) );
  OAI22XL U14708 ( .A0(n8174), .A1(n9036), .B0(n8170), .B1(n9034), .Y(n1912)
         );
  AOI221XL U14709 ( .A0(\xArray[13][46] ), .A1(n8179), .B0(\xArray[1][46] ), 
        .B1(n8177), .C0(n1903), .Y(n1902) );
  OAI22XL U14710 ( .A0(n8174), .A1(n9028), .B0(n8170), .B1(n9026), .Y(n1903)
         );
  AOI221XL U14711 ( .A0(\xArray[13][47] ), .A1(n8179), .B0(\xArray[1][47] ), 
        .B1(n8177), .C0(n1894), .Y(n1893) );
  OA22X1 U14712 ( .A0(n8319), .A1(n1362), .B0(n7713), .B1(n1601), .Y(n1892) );
  OAI22XL U14713 ( .A0(n8174), .A1(n9020), .B0(n8170), .B1(n9018), .Y(n1894)
         );
  MX4X1 U14714 ( .A(\bArray[8][48] ), .B(\bArray[9][48] ), .C(\bArray[10][48] ), .D(\bArray[11][48] ), .S0(n7200), .S1(n7213), .Y(n7137) );
  MX4X1 U14715 ( .A(\bArray[12][48] ), .B(\bArray[13][48] ), .C(
        \bArray[14][48] ), .D(\bArray[15][48] ), .S0(n7200), .S1(n7213), .Y(
        n7136) );
  MX4X1 U14716 ( .A(\bArray[4][48] ), .B(\bArray[5][48] ), .C(\bArray[6][48] ), 
        .D(\bArray[7][48] ), .S0(n7200), .S1(n7213), .Y(n7138) );
  OAI221X1 U14717 ( .A0(\xArray[7][52] ), .A1(n8285), .B0(\xArray[11][52] ), 
        .B1(n8225), .C0(n1034), .Y(n357) );
  OAI221X1 U14718 ( .A0(\xArray[7][53] ), .A1(n8296), .B0(\xArray[11][53] ), 
        .B1(n8225), .C0(n1029), .Y(n349) );
  OAI221X1 U14719 ( .A0(\xArray[7][54] ), .A1(n8296), .B0(\xArray[11][54] ), 
        .B1(n8225), .C0(n1024), .Y(n341) );
  OAI221X1 U14720 ( .A0(\xArray[4][53] ), .A1(n8280), .B0(\xArray[8][53] ), 
        .B1(n8226), .C0(n1846), .Y(n1336) );
  OAI221X1 U14721 ( .A0(\xArray[4][54] ), .A1(n8298), .B0(\xArray[8][54] ), 
        .B1(n8225), .C0(n1837), .Y(n1332) );
  OAI221X1 U14722 ( .A0(\xArray[4][55] ), .A1(n8287), .B0(\xArray[8][55] ), 
        .B1(n8232), .C0(n1828), .Y(n1328) );
  OAI221X1 U14723 ( .A0(\xArray[4][56] ), .A1(n8287), .B0(\xArray[8][56] ), 
        .B1(n8238), .C0(n1819), .Y(n1324) );
  OAI221X1 U14724 ( .A0(\xArray[8][52] ), .A1(n8297), .B0(\xArray[12][52] ), 
        .B1(n8225), .C0(n1033), .Y(n359) );
  OAI221X1 U14725 ( .A0(\xArray[8][53] ), .A1(n8293), .B0(\xArray[12][53] ), 
        .B1(n8225), .C0(n1028), .Y(n351) );
  OAI221X1 U14726 ( .A0(\xArray[8][54] ), .A1(n8296), .B0(\xArray[12][54] ), 
        .B1(n8225), .C0(n1023), .Y(n343) );
  OAI221X1 U14727 ( .A0(\xArray[6][53] ), .A1(n8279), .B0(\xArray[10][53] ), 
        .B1(n8233), .C0(n1339), .Y(n815) );
  OAI221X1 U14728 ( .A0(\xArray[6][54] ), .A1(n8279), .B0(\xArray[10][54] ), 
        .B1(n8233), .C0(n1335), .Y(n812) );
  OAI221X1 U14729 ( .A0(\xArray[5][53] ), .A1(n8286), .B0(\xArray[9][53] ), 
        .B1(n8227), .C0(n1584), .Y(n1027) );
  OAI221X1 U14730 ( .A0(\xArray[5][54] ), .A1(n8292), .B0(\xArray[9][54] ), 
        .B1(n8227), .C0(n1581), .Y(n1022) );
  OAI221X1 U14731 ( .A0(\xArray[5][55] ), .A1(n8286), .B0(\xArray[9][55] ), 
        .B1(n8225), .C0(n1578), .Y(n1017) );
  OAI221XL U14732 ( .A0(\xArray[9][51] ), .A1(n8281), .B0(\xArray[13][51] ), 
        .B1(n8238), .C0(n822), .Y(n366) );
  OAI221XL U14733 ( .A0(\xArray[9][52] ), .A1(n8281), .B0(\xArray[13][52] ), 
        .B1(n8232), .C0(n819), .Y(n358) );
  OAI221XL U14734 ( .A0(\xArray[2][51] ), .A1(n8286), .B0(\xArray[6][51] ), 
        .B1(n8233), .C0(n1861), .Y(n1589) );
  OAI222XL U14735 ( .A0(n429), .A1(n8338), .B0(n430), .B1(n8310), .C0(n431), 
        .C1(n7711), .Y(n424) );
  AOI221XL U14736 ( .A0(\xArray[14][43] ), .A1(n6573), .B0(\xArray[2][43] ), 
        .B1(n8360), .C0(n426), .Y(n425) );
  OAI22XL U14737 ( .A0(n8356), .A1(n9051), .B0(n8354), .B1(n9053), .Y(n426) );
  OAI222XL U14738 ( .A0(n437), .A1(n8338), .B0(n438), .B1(n8310), .C0(n439), 
        .C1(n7721), .Y(n432) );
  AOI221XL U14739 ( .A0(\xArray[14][42] ), .A1(n6573), .B0(\xArray[2][42] ), 
        .B1(n8360), .C0(n434), .Y(n433) );
  OAI22XL U14740 ( .A0(n8356), .A1(n9059), .B0(n8354), .B1(n9061), .Y(n434) );
  MX4X1 U14741 ( .A(n6928), .B(n6926), .C(n6927), .D(n6925), .S0(n7007), .S1(
        n8412), .Y(N25549) );
  MX4X1 U14742 ( .A(\bArray[8][51] ), .B(\bArray[9][51] ), .C(\bArray[10][51] ), .D(\bArray[11][51] ), .S0(n6989), .S1(n6994), .Y(n6926) );
  MX4X1 U14743 ( .A(\bArray[0][51] ), .B(\bArray[1][51] ), .C(\bArray[2][51] ), 
        .D(\bArray[3][51] ), .S0(n6989), .S1(n6994), .Y(n6928) );
  MX4X1 U14744 ( .A(\bArray[12][51] ), .B(\bArray[13][51] ), .C(
        \bArray[14][51] ), .D(\bArray[15][51] ), .S0(n6981), .S1(n6992), .Y(
        n6925) );
  MX4X1 U14745 ( .A(n6924), .B(n6922), .C(n6923), .D(n6921), .S0(n8411), .S1(
        n8412), .Y(N25550) );
  MX4X1 U14746 ( .A(\bArray[8][50] ), .B(\bArray[9][50] ), .C(\bArray[10][50] ), .D(\bArray[11][50] ), .S0(n6989), .S1(n7002), .Y(n6922) );
  MX4X1 U14747 ( .A(\bArray[0][50] ), .B(\bArray[1][50] ), .C(\bArray[2][50] ), 
        .D(\bArray[3][50] ), .S0(n6989), .S1(n7002), .Y(n6924) );
  MX4X1 U14748 ( .A(\bArray[12][50] ), .B(\bArray[13][50] ), .C(
        \bArray[14][50] ), .D(\bArray[15][50] ), .S0(n6989), .S1(n7002), .Y(
        n6921) );
  MX4X1 U14749 ( .A(n6920), .B(n6918), .C(n6919), .D(n6917), .S0(n8411), .S1(
        n8412), .Y(N25551) );
  MX4X1 U14750 ( .A(\bArray[8][49] ), .B(\bArray[9][49] ), .C(\bArray[10][49] ), .D(\bArray[11][49] ), .S0(n6981), .S1(n8413), .Y(n6918) );
  MX4X1 U14751 ( .A(\bArray[0][49] ), .B(\bArray[1][49] ), .C(\bArray[2][49] ), 
        .D(\bArray[3][49] ), .S0(n6977), .S1(n6992), .Y(n6920) );
  MX4X1 U14752 ( .A(\bArray[12][49] ), .B(\bArray[13][49] ), .C(
        \bArray[14][49] ), .D(\bArray[15][49] ), .S0(n8414), .S1(n7000), .Y(
        n6917) );
  MX4X1 U14753 ( .A(n6916), .B(n6914), .C(n6915), .D(n6913), .S0(n8411), .S1(
        n8412), .Y(N25552) );
  MX4X1 U14754 ( .A(\bArray[8][48] ), .B(\bArray[9][48] ), .C(\bArray[10][48] ), .D(\bArray[11][48] ), .S0(n8414), .S1(n7000), .Y(n6914) );
  MX4X1 U14755 ( .A(\bArray[0][48] ), .B(\bArray[1][48] ), .C(\bArray[2][48] ), 
        .D(\bArray[3][48] ), .S0(n8414), .S1(n7001), .Y(n6916) );
  MX4X1 U14756 ( .A(\bArray[12][48] ), .B(\bArray[13][48] ), .C(
        \bArray[14][48] ), .D(\bArray[15][48] ), .S0(n8414), .S1(n6993), .Y(
        n6913) );
  CLKINVX1 U14757 ( .A(\xArray[14][49] ), .Y(n9006) );
  CLKINVX1 U14758 ( .A(\xArray[14][50] ), .Y(n8998) );
  CLKINVX1 U14759 ( .A(\xArray[3][51] ), .Y(n8984) );
  MX4X1 U14760 ( .A(\bArray[4][51] ), .B(\bArray[5][51] ), .C(\bArray[6][51] ), 
        .D(\bArray[7][51] ), .S0(n6989), .S1(n6994), .Y(n6927) );
  MX4X1 U14761 ( .A(\bArray[4][50] ), .B(\bArray[5][50] ), .C(\bArray[6][50] ), 
        .D(\bArray[7][50] ), .S0(n6989), .S1(n7002), .Y(n6923) );
  MX4X1 U14762 ( .A(\bArray[4][49] ), .B(\bArray[5][49] ), .C(\bArray[6][49] ), 
        .D(\bArray[7][49] ), .S0(n6982), .S1(n7000), .Y(n6919) );
  MX4X1 U14763 ( .A(\bArray[4][48] ), .B(\bArray[5][48] ), .C(\bArray[6][48] ), 
        .D(\bArray[7][48] ), .S0(n8414), .S1(n7000), .Y(n6915) );
  MX4X1 U14764 ( .A(\bArray[0][48] ), .B(\bArray[1][48] ), .C(\bArray[2][48] ), 
        .D(\bArray[3][48] ), .S0(n7204), .S1(n7213), .Y(n7139) );
  OAI221X1 U14765 ( .A0(\xArray[3][53] ), .A1(n8286), .B0(\xArray[7][53] ), 
        .B1(n8233), .C0(n1845), .Y(n1338) );
  OAI221X1 U14766 ( .A0(\xArray[3][54] ), .A1(n8294), .B0(\xArray[7][54] ), 
        .B1(n8233), .C0(n1836), .Y(n1334) );
  OAI221X1 U14767 ( .A0(\xArray[3][55] ), .A1(n8287), .B0(\xArray[7][55] ), 
        .B1(n8237), .C0(n1827), .Y(n1330) );
  AOI221XL U14768 ( .A0(\xArray[13][48] ), .A1(n8179), .B0(\xArray[1][48] ), 
        .B1(n8177), .C0(n1885), .Y(n1884) );
  OA22X1 U14769 ( .A0(n8319), .A1(n1358), .B0(n7713), .B1(n1598), .Y(n1883) );
  OAI22XL U14770 ( .A0(n8174), .A1(n9012), .B0(n8170), .B1(n9010), .Y(n1885)
         );
  AOI221XL U14771 ( .A0(\xArray[13][49] ), .A1(n8179), .B0(\xArray[1][49] ), 
        .B1(n8177), .C0(n1876), .Y(n1875) );
  OA22X1 U14772 ( .A0(n8319), .A1(n1354), .B0(n7722), .B1(n1595), .Y(n1874) );
  OAI22XL U14773 ( .A0(n8174), .A1(n9004), .B0(n8170), .B1(n9002), .Y(n1876)
         );
  MX4X1 U14774 ( .A(\bArray[8][49] ), .B(\bArray[9][49] ), .C(\bArray[10][49] ), .D(\bArray[11][49] ), .S0(n7205), .S1(n7213), .Y(n7141) );
  MX4X1 U14775 ( .A(\bArray[12][49] ), .B(\bArray[13][49] ), .C(
        \bArray[14][49] ), .D(\bArray[15][49] ), .S0(n7205), .S1(n7213), .Y(
        n7140) );
  MX4X1 U14776 ( .A(\bArray[4][49] ), .B(\bArray[5][49] ), .C(\bArray[6][49] ), 
        .D(\bArray[7][49] ), .S0(n7200), .S1(n7213), .Y(n7142) );
  MX4X1 U14777 ( .A(\bArray[8][50] ), .B(\bArray[9][50] ), .C(\bArray[10][50] ), .D(\bArray[11][50] ), .S0(n7202), .S1(n7213), .Y(n7145) );
  MX4X1 U14778 ( .A(\bArray[12][50] ), .B(\bArray[13][50] ), .C(
        \bArray[14][50] ), .D(\bArray[15][50] ), .S0(n7200), .S1(n7213), .Y(
        n7144) );
  MX4X1 U14779 ( .A(\bArray[4][50] ), .B(\bArray[5][50] ), .C(\bArray[6][50] ), 
        .D(\bArray[7][50] ), .S0(n7202), .S1(n7214), .Y(n7146) );
  MX4X1 U14780 ( .A(\bArray[8][51] ), .B(\bArray[9][51] ), .C(\bArray[10][51] ), .D(\bArray[11][51] ), .S0(n7201), .S1(N1762), .Y(n7149) );
  MX4X1 U14781 ( .A(\bArray[12][51] ), .B(\bArray[13][51] ), .C(
        \bArray[14][51] ), .D(\bArray[15][51] ), .S0(n7202), .S1(N1762), .Y(
        n7148) );
  MX4X1 U14782 ( .A(\bArray[4][51] ), .B(\bArray[5][51] ), .C(\bArray[6][51] ), 
        .D(\bArray[7][51] ), .S0(n7211), .S1(N1762), .Y(n7150) );
  OAI221X1 U14783 ( .A0(\xArray[7][55] ), .A1(n8296), .B0(\xArray[11][55] ), 
        .B1(n8225), .C0(n1019), .Y(n333) );
  OAI221X1 U14784 ( .A0(\xArray[7][56] ), .A1(n8289), .B0(\xArray[11][56] ), 
        .B1(n8235), .C0(n1014), .Y(n325) );
  AOI2BB2X1 U14785 ( .B0(n8944), .B1(n8209), .A0N(\xArray[15][56] ), .A1N(
        n8259), .Y(n1014) );
  OAI221X1 U14786 ( .A0(\xArray[4][57] ), .A1(n8287), .B0(\xArray[8][57] ), 
        .B1(n8236), .C0(n1810), .Y(n1320) );
  OAI221X1 U14787 ( .A0(\xArray[8][55] ), .A1(n8296), .B0(\xArray[12][55] ), 
        .B1(n8225), .C0(n1018), .Y(n335) );
  OAI221X1 U14788 ( .A0(\xArray[8][56] ), .A1(n8289), .B0(\xArray[12][56] ), 
        .B1(n8235), .C0(n1013), .Y(n327) );
  OAI221X1 U14789 ( .A0(\xArray[6][55] ), .A1(n8279), .B0(\xArray[10][55] ), 
        .B1(n8237), .C0(n1331), .Y(n809) );
  OAI221X1 U14790 ( .A0(\xArray[6][56] ), .A1(n8279), .B0(\xArray[10][56] ), 
        .B1(n8237), .C0(n1327), .Y(n806) );
  OAI221X1 U14791 ( .A0(\xArray[6][57] ), .A1(n8279), .B0(\xArray[10][57] ), 
        .B1(n8243), .C0(n1323), .Y(n803) );
  OAI221X1 U14792 ( .A0(\xArray[5][56] ), .A1(n8295), .B0(\xArray[9][56] ), 
        .B1(n8227), .C0(n1575), .Y(n1012) );
  OAI221X1 U14793 ( .A0(\xArray[5][57] ), .A1(n8292), .B0(\xArray[9][57] ), 
        .B1(n8227), .C0(n1572), .Y(n1007) );
  OAI221XL U14794 ( .A0(\xArray[9][53] ), .A1(n8281), .B0(\xArray[13][53] ), 
        .B1(n8241), .C0(n816), .Y(n350) );
  OAI221XL U14795 ( .A0(\xArray[9][54] ), .A1(n8289), .B0(\xArray[13][54] ), 
        .B1(n8238), .C0(n813), .Y(n342) );
  OAI221XL U14796 ( .A0(\xArray[2][52] ), .A1(n8286), .B0(\xArray[6][52] ), 
        .B1(n8233), .C0(n1852), .Y(n1586) );
  OAI221XL U14797 ( .A0(\xArray[2][53] ), .A1(n8278), .B0(\xArray[6][53] ), 
        .B1(n8233), .C0(n1843), .Y(n1583) );
  OAI222XL U14798 ( .A0(n413), .A1(n8338), .B0(n414), .B1(n8310), .C0(n415), 
        .C1(n7707), .Y(n408) );
  AOI221XL U14799 ( .A0(\xArray[14][45] ), .A1(n6573), .B0(\xArray[2][45] ), 
        .B1(n8360), .C0(n410), .Y(n409) );
  OAI22XL U14800 ( .A0(n8356), .A1(n9035), .B0(n8354), .B1(n9037), .Y(n410) );
  OAI222XL U14801 ( .A0(n421), .A1(n8338), .B0(n422), .B1(n8310), .C0(n423), 
        .C1(n7707), .Y(n416) );
  AOI221XL U14802 ( .A0(\xArray[14][44] ), .A1(n6573), .B0(\xArray[2][44] ), 
        .B1(n8360), .C0(n418), .Y(n417) );
  OAI22XL U14803 ( .A0(n8356), .A1(n9043), .B0(n8354), .B1(n9045), .Y(n418) );
  CLKINVX1 U14804 ( .A(\xArray[14][51] ), .Y(n8990) );
  CLKINVX1 U14805 ( .A(\xArray[14][52] ), .Y(n8982) );
  CLKINVX1 U14806 ( .A(\xArray[5][44] ), .Y(n9042) );
  CLKINVX1 U14807 ( .A(\xArray[5][45] ), .Y(n9034) );
  CLKINVX1 U14808 ( .A(\xArray[5][46] ), .Y(n9026) );
  CLKINVX1 U14809 ( .A(\xArray[5][47] ), .Y(n9018) );
  CLKINVX1 U14810 ( .A(\xArray[3][52] ), .Y(n8976) );
  CLKINVX1 U14811 ( .A(\xArray[3][53] ), .Y(n8968) );
  CLKINVX1 U14812 ( .A(\xArray[3][54] ), .Y(n8960) );
  MX4X1 U14813 ( .A(\bArray[0][49] ), .B(\bArray[1][49] ), .C(\bArray[2][49] ), 
        .D(\bArray[3][49] ), .S0(n7200), .S1(n7213), .Y(n7143) );
  MX4X1 U14814 ( .A(\bArray[0][50] ), .B(\bArray[1][50] ), .C(\bArray[2][50] ), 
        .D(\bArray[3][50] ), .S0(n7200), .S1(n7213), .Y(n7147) );
  MX4X1 U14815 ( .A(\bArray[0][51] ), .B(\bArray[1][51] ), .C(\bArray[2][51] ), 
        .D(\bArray[3][51] ), .S0(n7209), .S1(N1762), .Y(n7151) );
  CLKINVX1 U14816 ( .A(\xArray[9][44] ), .Y(n9044) );
  CLKINVX1 U14817 ( .A(\xArray[9][45] ), .Y(n9036) );
  CLKINVX1 U14818 ( .A(\xArray[9][46] ), .Y(n9028) );
  CLKINVX1 U14819 ( .A(\xArray[9][47] ), .Y(n9020) );
  OAI221X1 U14820 ( .A0(\xArray[3][56] ), .A1(n8287), .B0(\xArray[7][56] ), 
        .B1(n8235), .C0(n1818), .Y(n1326) );
  OAI221X1 U14821 ( .A0(\xArray[3][57] ), .A1(n8287), .B0(\xArray[7][57] ), 
        .B1(n8241), .C0(n1809), .Y(n1322) );
  CLKINVX1 U14822 ( .A(\xArray[6][43] ), .Y(n9051) );
  CLKINVX1 U14823 ( .A(\xArray[6][42] ), .Y(n9059) );
  CLKINVX1 U14824 ( .A(\xArray[10][43] ), .Y(n9053) );
  CLKINVX1 U14825 ( .A(\xArray[10][42] ), .Y(n9061) );
  AOI221XL U14826 ( .A0(\xArray[13][50] ), .A1(n8179), .B0(\xArray[1][50] ), 
        .B1(n8177), .C0(n1867), .Y(n1866) );
  OA22X1 U14827 ( .A0(n8319), .A1(n1350), .B0(n7730), .B1(n1592), .Y(n1865) );
  OAI22XL U14828 ( .A0(n8174), .A1(n8996), .B0(n8170), .B1(n8994), .Y(n1867)
         );
  AOI221XL U14829 ( .A0(\xArray[13][51] ), .A1(n8179), .B0(\xArray[1][51] ), 
        .B1(n8177), .C0(n1858), .Y(n1857) );
  OAI22XL U14830 ( .A0(n8174), .A1(n8988), .B0(n8170), .B1(n8986), .Y(n1858)
         );
  MX4X1 U14831 ( .A(\bArray[8][52] ), .B(\bArray[9][52] ), .C(\bArray[10][52] ), .D(\bArray[11][52] ), .S0(n7211), .S1(n7215), .Y(n7153) );
  MX4X1 U14832 ( .A(\bArray[12][52] ), .B(\bArray[13][52] ), .C(
        \bArray[14][52] ), .D(\bArray[15][52] ), .S0(n7211), .S1(n7215), .Y(
        n7152) );
  MX4X1 U14833 ( .A(\bArray[4][52] ), .B(\bArray[5][52] ), .C(\bArray[6][52] ), 
        .D(\bArray[7][52] ), .S0(n7211), .S1(n7215), .Y(n7154) );
  OAI221X1 U14834 ( .A0(\xArray[7][57] ), .A1(n8289), .B0(\xArray[11][57] ), 
        .B1(n8235), .C0(n1009), .Y(n317) );
  AOI2BB2X1 U14835 ( .B0(n8936), .B1(n8208), .A0N(\xArray[15][57] ), .A1N(
        n8259), .Y(n1009) );
  OAI221X1 U14836 ( .A0(\xArray[7][58] ), .A1(n8289), .B0(\xArray[11][58] ), 
        .B1(n8235), .C0(n1004), .Y(n309) );
  AOI2BB2X1 U14837 ( .B0(n8928), .B1(n8208), .A0N(\xArray[15][58] ), .A1N(
        n8259), .Y(n1004) );
  OAI221X1 U14838 ( .A0(\xArray[4][58] ), .A1(n8287), .B0(\xArray[8][58] ), 
        .B1(n8226), .C0(n1801), .Y(n1316) );
  OAI221X1 U14839 ( .A0(\xArray[4][59] ), .A1(n8287), .B0(\xArray[8][59] ), 
        .B1(n8229), .C0(n1792), .Y(n1312) );
  OAI221X1 U14840 ( .A0(\xArray[4][60] ), .A1(n8280), .B0(\xArray[8][60] ), 
        .B1(n8226), .C0(n1783), .Y(n1308) );
  OAI221X1 U14841 ( .A0(\xArray[8][57] ), .A1(n8289), .B0(\xArray[12][57] ), 
        .B1(n8235), .C0(n1008), .Y(n319) );
  OAI221X1 U14842 ( .A0(\xArray[8][58] ), .A1(n8289), .B0(\xArray[12][58] ), 
        .B1(n8235), .C0(n1003), .Y(n311) );
  OAI221X1 U14843 ( .A0(\xArray[6][58] ), .A1(n8279), .B0(\xArray[10][58] ), 
        .B1(n8231), .C0(n1319), .Y(n800) );
  OAI221X1 U14844 ( .A0(\xArray[6][59] ), .A1(n8279), .B0(\xArray[10][59] ), 
        .B1(n8231), .C0(n1315), .Y(n797) );
  OAI221X1 U14845 ( .A0(\xArray[5][58] ), .A1(n8286), .B0(\xArray[9][58] ), 
        .B1(n8227), .C0(n1569), .Y(n1002) );
  OAI221X1 U14846 ( .A0(\xArray[5][59] ), .A1(n8283), .B0(\xArray[9][59] ), 
        .B1(n8229), .C0(n1566), .Y(n997) );
  OA22X1 U14847 ( .A0(\xArray[1][59] ), .A1(n8199), .B0(\xArray[13][59] ), 
        .B1(n8267), .Y(n1566) );
  OAI221XL U14848 ( .A0(\xArray[9][55] ), .A1(n8292), .B0(\xArray[13][55] ), 
        .B1(n8238), .C0(n810), .Y(n334) );
  OA22X1 U14849 ( .A0(\xArray[5][55] ), .A1(n8194), .B0(\xArray[1][55] ), .B1(
        n8254), .Y(n810) );
  OAI221XL U14850 ( .A0(\xArray[9][56] ), .A1(n8292), .B0(\xArray[13][56] ), 
        .B1(n8238), .C0(n807), .Y(n326) );
  OA22X1 U14851 ( .A0(\xArray[5][56] ), .A1(n8194), .B0(\xArray[1][56] ), .B1(
        n8254), .Y(n807) );
  OAI221XL U14852 ( .A0(\xArray[2][54] ), .A1(n8298), .B0(\xArray[6][54] ), 
        .B1(n8233), .C0(n1834), .Y(n1580) );
  OAI221XL U14853 ( .A0(\xArray[2][55] ), .A1(n8298), .B0(\xArray[6][55] ), 
        .B1(n8233), .C0(n1825), .Y(n1577) );
  OAI221XL U14854 ( .A0(\xArray[2][56] ), .A1(n8287), .B0(\xArray[6][56] ), 
        .B1(n8241), .C0(n1816), .Y(n1574) );
  OAI222XL U14855 ( .A0(n397), .A1(n8338), .B0(n398), .B1(n8310), .C0(n399), 
        .C1(n7713), .Y(n392) );
  AOI221XL U14856 ( .A0(\xArray[14][47] ), .A1(n6573), .B0(\xArray[2][47] ), 
        .B1(n8360), .C0(n394), .Y(n393) );
  OAI22XL U14857 ( .A0(n8356), .A1(n9019), .B0(n8354), .B1(n9021), .Y(n394) );
  OAI222XL U14858 ( .A0(n405), .A1(n8338), .B0(n406), .B1(n8310), .C0(n407), 
        .C1(n7740), .Y(n400) );
  AOI221XL U14859 ( .A0(\xArray[14][46] ), .A1(n6573), .B0(\xArray[2][46] ), 
        .B1(n8360), .C0(n402), .Y(n401) );
  OAI22XL U14860 ( .A0(n8356), .A1(n9027), .B0(n8354), .B1(n9029), .Y(n402) );
  MX4X1 U14861 ( .A(n6944), .B(n6942), .C(n6943), .D(n6941), .S0(n7007), .S1(
        n7004), .Y(N25545) );
  MX4X1 U14862 ( .A(\bArray[8][55] ), .B(\bArray[9][55] ), .C(\bArray[10][55] ), .D(\bArray[11][55] ), .S0(N1757), .S1(n6993), .Y(n6942) );
  MX4X1 U14863 ( .A(\bArray[0][55] ), .B(\bArray[1][55] ), .C(\bArray[2][55] ), 
        .D(\bArray[3][55] ), .S0(N1757), .S1(n6993), .Y(n6944) );
  MX4X1 U14864 ( .A(\bArray[12][55] ), .B(\bArray[13][55] ), .C(
        \bArray[14][55] ), .D(\bArray[15][55] ), .S0(n8414), .S1(n6993), .Y(
        n6941) );
  MX4X1 U14865 ( .A(n6940), .B(n6938), .C(n6939), .D(n6937), .S0(n7007), .S1(
        n7004), .Y(N25546) );
  MX4X1 U14866 ( .A(\bArray[8][54] ), .B(\bArray[9][54] ), .C(\bArray[10][54] ), .D(\bArray[11][54] ), .S0(n6983), .S1(n6993), .Y(n6938) );
  MX4X1 U14867 ( .A(\bArray[0][54] ), .B(\bArray[1][54] ), .C(\bArray[2][54] ), 
        .D(\bArray[3][54] ), .S0(n6981), .S1(n6993), .Y(n6940) );
  MX4X1 U14868 ( .A(\bArray[12][54] ), .B(\bArray[13][54] ), .C(
        \bArray[14][54] ), .D(\bArray[15][54] ), .S0(n6982), .S1(n7001), .Y(
        n6937) );
  MX4X1 U14869 ( .A(n6936), .B(n6934), .C(n6935), .D(n6933), .S0(n7007), .S1(
        n8412), .Y(N25547) );
  MX4X1 U14870 ( .A(\bArray[8][53] ), .B(\bArray[9][53] ), .C(\bArray[10][53] ), .D(\bArray[11][53] ), .S0(n6977), .S1(n6995), .Y(n6934) );
  MX4X1 U14871 ( .A(\bArray[0][53] ), .B(\bArray[1][53] ), .C(\bArray[2][53] ), 
        .D(\bArray[3][53] ), .S0(n6982), .S1(n6995), .Y(n6936) );
  MX4X1 U14872 ( .A(\bArray[12][53] ), .B(\bArray[13][53] ), .C(
        \bArray[14][53] ), .D(\bArray[15][53] ), .S0(n6989), .S1(n6995), .Y(
        n6933) );
  MX4X1 U14873 ( .A(n6932), .B(n6930), .C(n6931), .D(n6929), .S0(n7007), .S1(
        n8412), .Y(N25548) );
  MX4X1 U14874 ( .A(\bArray[8][52] ), .B(\bArray[9][52] ), .C(\bArray[10][52] ), .D(\bArray[11][52] ), .S0(n6989), .S1(n6994), .Y(n6930) );
  MX4X1 U14875 ( .A(\bArray[0][52] ), .B(\bArray[1][52] ), .C(\bArray[2][52] ), 
        .D(\bArray[3][52] ), .S0(n6989), .S1(n6995), .Y(n6932) );
  MX4X1 U14876 ( .A(\bArray[12][52] ), .B(\bArray[13][52] ), .C(
        \bArray[14][52] ), .D(\bArray[15][52] ), .S0(n6989), .S1(n6994), .Y(
        n6929) );
  CLKINVX1 U14877 ( .A(\xArray[14][53] ), .Y(n8974) );
  CLKINVX1 U14878 ( .A(\xArray[14][54] ), .Y(n8966) );
  CLKINVX1 U14879 ( .A(\xArray[3][55] ), .Y(n8952) );
  CLKINVX1 U14880 ( .A(\xArray[3][56] ), .Y(n8944) );
  MX4X1 U14881 ( .A(\bArray[4][55] ), .B(\bArray[5][55] ), .C(\bArray[6][55] ), 
        .D(\bArray[7][55] ), .S0(N1757), .S1(n6993), .Y(n6943) );
  MX4X1 U14882 ( .A(\bArray[4][54] ), .B(\bArray[5][54] ), .C(\bArray[6][54] ), 
        .D(\bArray[7][54] ), .S0(n6990), .S1(n6993), .Y(n6939) );
  MX4X1 U14883 ( .A(\bArray[4][53] ), .B(\bArray[5][53] ), .C(\bArray[6][53] ), 
        .D(\bArray[7][53] ), .S0(n6989), .S1(n6995), .Y(n6935) );
  MX4X1 U14884 ( .A(\bArray[4][52] ), .B(\bArray[5][52] ), .C(\bArray[6][52] ), 
        .D(\bArray[7][52] ), .S0(n6989), .S1(n6994), .Y(n6931) );
  MX4X1 U14885 ( .A(\bArray[0][52] ), .B(\bArray[1][52] ), .C(\bArray[2][52] ), 
        .D(\bArray[3][52] ), .S0(n7211), .S1(n7215), .Y(n7155) );
  OAI221X1 U14886 ( .A0(\xArray[3][58] ), .A1(n8287), .B0(\xArray[7][58] ), 
        .B1(n8226), .C0(n1800), .Y(n1318) );
  OAI221X1 U14887 ( .A0(\xArray[3][59] ), .A1(n8287), .B0(\xArray[7][59] ), 
        .B1(n8226), .C0(n1791), .Y(n1314) );
  AOI221XL U14888 ( .A0(\xArray[13][52] ), .A1(n8179), .B0(\xArray[1][52] ), 
        .B1(n8177), .C0(n1849), .Y(n1848) );
  OAI22XL U14889 ( .A0(n8173), .A1(n8980), .B0(n8170), .B1(n8978), .Y(n1849)
         );
  AOI221XL U14890 ( .A0(\xArray[13][53] ), .A1(n8179), .B0(\xArray[1][53] ), 
        .B1(n8176), .C0(n1840), .Y(n1839) );
  OAI22XL U14891 ( .A0(n8173), .A1(n8972), .B0(n8170), .B1(n8970), .Y(n1840)
         );
  MX4X1 U14892 ( .A(\bArray[8][53] ), .B(\bArray[9][53] ), .C(\bArray[10][53] ), .D(\bArray[11][53] ), .S0(n7201), .S1(n7214), .Y(n7157) );
  MX4X1 U14893 ( .A(\bArray[12][53] ), .B(\bArray[13][53] ), .C(
        \bArray[14][53] ), .D(\bArray[15][53] ), .S0(n7211), .S1(n7221), .Y(
        n7156) );
  MX4X1 U14894 ( .A(\bArray[4][53] ), .B(\bArray[5][53] ), .C(\bArray[6][53] ), 
        .D(\bArray[7][53] ), .S0(n7201), .S1(n7214), .Y(n7158) );
  MX4X1 U14895 ( .A(\bArray[8][54] ), .B(\bArray[9][54] ), .C(\bArray[10][54] ), .D(\bArray[11][54] ), .S0(n7207), .S1(n7222), .Y(n7161) );
  MX4X1 U14896 ( .A(\bArray[12][54] ), .B(\bArray[13][54] ), .C(
        \bArray[14][54] ), .D(\bArray[15][54] ), .S0(n7201), .S1(n8409), .Y(
        n7160) );
  MX4X1 U14897 ( .A(\bArray[4][54] ), .B(\bArray[5][54] ), .C(\bArray[6][54] ), 
        .D(\bArray[7][54] ), .S0(n7207), .S1(n7222), .Y(n7162) );
  MX4X1 U14898 ( .A(\bArray[8][55] ), .B(\bArray[9][55] ), .C(\bArray[10][55] ), .D(\bArray[11][55] ), .S0(n7207), .S1(n7212), .Y(n7165) );
  MX4X1 U14899 ( .A(\bArray[12][55] ), .B(\bArray[13][55] ), .C(
        \bArray[14][55] ), .D(\bArray[15][55] ), .S0(n7207), .S1(n7212), .Y(
        n7164) );
  MX4X1 U14900 ( .A(\bArray[4][55] ), .B(\bArray[5][55] ), .C(\bArray[6][55] ), 
        .D(\bArray[7][55] ), .S0(n7207), .S1(n7212), .Y(n7166) );
  OAI221X1 U14901 ( .A0(\xArray[7][60] ), .A1(n8289), .B0(\xArray[11][60] ), 
        .B1(n8235), .C0(n994), .Y(n293) );
  OAI221X1 U14902 ( .A0(\xArray[7][59] ), .A1(n8289), .B0(\xArray[11][59] ), 
        .B1(n8235), .C0(n999), .Y(n301) );
  OAI221X1 U14903 ( .A0(\xArray[8][59] ), .A1(n8289), .B0(\xArray[12][59] ), 
        .B1(n8235), .C0(n998), .Y(n303) );
  OAI221X1 U14904 ( .A0(\xArray[3][60] ), .A1(n8280), .B0(\xArray[7][60] ), 
        .B1(n8226), .C0(n1782), .Y(n1310) );
  OAI221X1 U14905 ( .A0(\xArray[6][60] ), .A1(n8279), .B0(\xArray[10][60] ), 
        .B1(n8239), .C0(n1311), .Y(n794) );
  OAI221X1 U14906 ( .A0(\xArray[5][60] ), .A1(n8283), .B0(\xArray[9][60] ), 
        .B1(n8229), .C0(n1563), .Y(n992) );
  OA22X1 U14907 ( .A0(\xArray[1][60] ), .A1(n8199), .B0(\xArray[13][60] ), 
        .B1(n8267), .Y(n1563) );
  OAI221XL U14908 ( .A0(\xArray[9][57] ), .A1(n8292), .B0(\xArray[13][57] ), 
        .B1(n8238), .C0(n804), .Y(n318) );
  OA22X1 U14909 ( .A0(\xArray[5][57] ), .A1(n8194), .B0(\xArray[1][57] ), .B1(
        n8254), .Y(n804) );
  OAI221XL U14910 ( .A0(\xArray[2][57] ), .A1(n8287), .B0(\xArray[6][57] ), 
        .B1(n8232), .C0(n1807), .Y(n1571) );
  OAI221XL U14911 ( .A0(\xArray[2][58] ), .A1(n8287), .B0(\xArray[6][58] ), 
        .B1(n8236), .C0(n1798), .Y(n1568) );
  OAI222XL U14912 ( .A0(n381), .A1(n8337), .B0(n382), .B1(n8307), .C0(n383), 
        .C1(n7730), .Y(n376) );
  AOI221XL U14913 ( .A0(\xArray[14][49] ), .A1(n6573), .B0(\xArray[2][49] ), 
        .B1(n8360), .C0(n378), .Y(n377) );
  OAI22XL U14914 ( .A0(n8356), .A1(n9003), .B0(n8354), .B1(n9005), .Y(n378) );
  OAI222XL U14915 ( .A0(n389), .A1(n8337), .B0(n390), .B1(n8306), .C0(n391), 
        .C1(n7713), .Y(n384) );
  AOI221XL U14916 ( .A0(\xArray[14][48] ), .A1(n6573), .B0(\xArray[2][48] ), 
        .B1(n8360), .C0(n386), .Y(n385) );
  OAI22XL U14917 ( .A0(n8356), .A1(n9011), .B0(n8354), .B1(n9013), .Y(n386) );
  CLKINVX1 U14918 ( .A(\xArray[14][55] ), .Y(n8958) );
  CLKINVX1 U14919 ( .A(\xArray[14][56] ), .Y(n8950) );
  CLKINVX1 U14920 ( .A(\xArray[5][48] ), .Y(n9010) );
  CLKINVX1 U14921 ( .A(\xArray[5][49] ), .Y(n9002) );
  CLKINVX1 U14922 ( .A(\xArray[5][50] ), .Y(n8994) );
  CLKINVX1 U14923 ( .A(\xArray[5][51] ), .Y(n8986) );
  CLKINVX1 U14924 ( .A(\xArray[3][57] ), .Y(n8936) );
  CLKINVX1 U14925 ( .A(\xArray[3][58] ), .Y(n8928) );
  MX4X1 U14926 ( .A(\bArray[0][53] ), .B(\bArray[1][53] ), .C(\bArray[2][53] ), 
        .D(\bArray[3][53] ), .S0(n7211), .S1(n7214), .Y(n7159) );
  MX4X1 U14927 ( .A(\bArray[0][54] ), .B(\bArray[1][54] ), .C(\bArray[2][54] ), 
        .D(\bArray[3][54] ), .S0(n7207), .S1(n7213), .Y(n7163) );
  MX4X1 U14928 ( .A(\bArray[0][55] ), .B(\bArray[1][55] ), .C(\bArray[2][55] ), 
        .D(\bArray[3][55] ), .S0(n7207), .S1(n7222), .Y(n7167) );
  CLKINVX1 U14929 ( .A(\xArray[9][48] ), .Y(n9012) );
  CLKINVX1 U14930 ( .A(\xArray[9][49] ), .Y(n9004) );
  CLKINVX1 U14931 ( .A(\xArray[9][50] ), .Y(n8996) );
  CLKINVX1 U14932 ( .A(\xArray[9][51] ), .Y(n8988) );
  CLKINVX1 U14933 ( .A(\xArray[6][47] ), .Y(n9019) );
  CLKINVX1 U14934 ( .A(\xArray[6][46] ), .Y(n9027) );
  CLKINVX1 U14935 ( .A(\xArray[6][45] ), .Y(n9035) );
  CLKINVX1 U14936 ( .A(\xArray[6][44] ), .Y(n9043) );
  CLKINVX1 U14937 ( .A(\xArray[10][47] ), .Y(n9021) );
  CLKINVX1 U14938 ( .A(\xArray[10][46] ), .Y(n9029) );
  CLKINVX1 U14939 ( .A(\xArray[10][45] ), .Y(n9037) );
  CLKINVX1 U14940 ( .A(\xArray[10][44] ), .Y(n9045) );
  AOI221XL U14941 ( .A0(\xArray[13][54] ), .A1(n8179), .B0(\xArray[1][54] ), 
        .B1(n8176), .C0(n1831), .Y(n1830) );
  OAI22XL U14942 ( .A0(n8173), .A1(n8964), .B0(n8172), .B1(n8962), .Y(n1831)
         );
  AOI221XL U14943 ( .A0(\xArray[13][55] ), .A1(n8179), .B0(\xArray[1][55] ), 
        .B1(n1747), .C0(n1822), .Y(n1821) );
  OAI22XL U14944 ( .A0(n8173), .A1(n8956), .B0(n8172), .B1(n8954), .Y(n1822)
         );
  MX4X1 U14945 ( .A(\bArray[8][56] ), .B(\bArray[9][56] ), .C(\bArray[10][56] ), .D(\bArray[11][56] ), .S0(n7203), .S1(n7212), .Y(n7169) );
  MX4X1 U14946 ( .A(\bArray[12][56] ), .B(\bArray[13][56] ), .C(
        \bArray[14][56] ), .D(\bArray[15][56] ), .S0(n7203), .S1(n7212), .Y(
        n7168) );
  MX4X1 U14947 ( .A(\bArray[4][56] ), .B(\bArray[5][56] ), .C(\bArray[6][56] ), 
        .D(\bArray[7][56] ), .S0(n7203), .S1(n7213), .Y(n7170) );
  OAI221X1 U14948 ( .A0(\xArray[7][61] ), .A1(n8289), .B0(\xArray[11][61] ), 
        .B1(n8235), .C0(n989), .Y(n285) );
  OAI221X1 U14949 ( .A0(\xArray[4][61] ), .A1(n8280), .B0(\xArray[8][61] ), 
        .B1(n8226), .C0(n1774), .Y(n1304) );
  OAI221X1 U14950 ( .A0(\xArray[8][61] ), .A1(n8289), .B0(\xArray[12][61] ), 
        .B1(n8235), .C0(n988), .Y(n287) );
  OAI221X1 U14951 ( .A0(\xArray[6][61] ), .A1(n8279), .B0(\xArray[10][61] ), 
        .B1(n8242), .C0(n1307), .Y(n791) );
  OAI221X1 U14952 ( .A0(\xArray[3][61] ), .A1(n8280), .B0(\xArray[7][61] ), 
        .B1(n8226), .C0(n1773), .Y(n1306) );
  OAI221X1 U14953 ( .A0(\xArray[5][61] ), .A1(n8283), .B0(\xArray[9][61] ), 
        .B1(n8229), .C0(n1560), .Y(n987) );
  OA22X1 U14954 ( .A0(\xArray[1][61] ), .A1(n8198), .B0(\xArray[13][61] ), 
        .B1(n8267), .Y(n1560) );
  OAI221XL U14955 ( .A0(\xArray[9][58] ), .A1(n8292), .B0(\xArray[13][58] ), 
        .B1(n8238), .C0(n801), .Y(n310) );
  OA22X1 U14956 ( .A0(\xArray[5][58] ), .A1(n8198), .B0(\xArray[1][58] ), .B1(
        n8258), .Y(n801) );
  OAI221XL U14957 ( .A0(\xArray[9][59] ), .A1(n8292), .B0(\xArray[13][59] ), 
        .B1(n8238), .C0(n798), .Y(n302) );
  OA22X1 U14958 ( .A0(\xArray[5][59] ), .A1(n8198), .B0(\xArray[1][59] ), .B1(
        n8254), .Y(n798) );
  OAI221XL U14959 ( .A0(\xArray[2][59] ), .A1(n8287), .B0(\xArray[6][59] ), 
        .B1(n8236), .C0(n1789), .Y(n1565) );
  OAI222XL U14960 ( .A0(n365), .A1(n8337), .B0(n366), .B1(n268), .C0(n367), 
        .C1(n7713), .Y(n360) );
  AOI221XL U14961 ( .A0(\xArray[14][51] ), .A1(n6573), .B0(\xArray[2][51] ), 
        .B1(n8360), .C0(n362), .Y(n361) );
  OAI22XL U14962 ( .A0(n8356), .A1(n8987), .B0(n8354), .B1(n8989), .Y(n362) );
  OAI222XL U14963 ( .A0(n373), .A1(n8337), .B0(n374), .B1(n8307), .C0(n375), 
        .C1(n7733), .Y(n368) );
  AOI221XL U14964 ( .A0(\xArray[14][50] ), .A1(n6573), .B0(\xArray[2][50] ), 
        .B1(n8360), .C0(n370), .Y(n369) );
  OAI22XL U14965 ( .A0(n8356), .A1(n8995), .B0(n8354), .B1(n8997), .Y(n370) );
  MX4X1 U14966 ( .A(n6960), .B(n6958), .C(n6959), .D(n6957), .S0(n7007), .S1(
        n8412), .Y(N25541) );
  MX4X1 U14967 ( .A(\bArray[8][59] ), .B(\bArray[9][59] ), .C(\bArray[10][59] ), .D(\bArray[11][59] ), .S0(n6978), .S1(n7002), .Y(n6958) );
  MX4X1 U14968 ( .A(\bArray[0][59] ), .B(\bArray[1][59] ), .C(\bArray[2][59] ), 
        .D(\bArray[3][59] ), .S0(n6985), .S1(n7002), .Y(n6960) );
  MX4X1 U14969 ( .A(\bArray[12][59] ), .B(\bArray[13][59] ), .C(
        \bArray[14][59] ), .D(\bArray[15][59] ), .S0(n6985), .S1(n7002), .Y(
        n6957) );
  MX4X1 U14970 ( .A(n6956), .B(n6954), .C(n6955), .D(n6953), .S0(n7007), .S1(
        n7004), .Y(N25542) );
  MX4X1 U14971 ( .A(\bArray[8][58] ), .B(\bArray[9][58] ), .C(\bArray[10][58] ), .D(\bArray[11][58] ), .S0(n6990), .S1(n6994), .Y(n6954) );
  MX4X1 U14972 ( .A(\bArray[0][58] ), .B(\bArray[1][58] ), .C(\bArray[2][58] ), 
        .D(\bArray[3][58] ), .S0(n6990), .S1(n6994), .Y(n6956) );
  MX4X1 U14973 ( .A(\bArray[12][58] ), .B(\bArray[13][58] ), .C(
        \bArray[14][58] ), .D(\bArray[15][58] ), .S0(n6990), .S1(n6994), .Y(
        n6953) );
  MX4X1 U14974 ( .A(n6952), .B(n6950), .C(n6951), .D(n6949), .S0(n7007), .S1(
        n7004), .Y(N25543) );
  MX4X1 U14975 ( .A(\bArray[8][57] ), .B(\bArray[9][57] ), .C(\bArray[10][57] ), .D(\bArray[11][57] ), .S0(n6990), .S1(n7001), .Y(n6950) );
  MX4X1 U14976 ( .A(\bArray[0][57] ), .B(\bArray[1][57] ), .C(\bArray[2][57] ), 
        .D(\bArray[3][57] ), .S0(n6990), .S1(n6994), .Y(n6952) );
  MX4X1 U14977 ( .A(\bArray[12][57] ), .B(\bArray[13][57] ), .C(
        \bArray[14][57] ), .D(\bArray[15][57] ), .S0(n8414), .S1(n7000), .Y(
        n6949) );
  MX4X1 U14978 ( .A(n6948), .B(n6946), .C(n6947), .D(n6945), .S0(n7007), .S1(
        n7003), .Y(N25544) );
  MX4X1 U14979 ( .A(\bArray[8][56] ), .B(\bArray[9][56] ), .C(\bArray[10][56] ), .D(\bArray[11][56] ), .S0(n8414), .S1(n7001), .Y(n6946) );
  MX4X1 U14980 ( .A(\bArray[0][56] ), .B(\bArray[1][56] ), .C(\bArray[2][56] ), 
        .D(\bArray[3][56] ), .S0(n8414), .S1(n6993), .Y(n6948) );
  MX4X1 U14981 ( .A(\bArray[12][56] ), .B(\bArray[13][56] ), .C(
        \bArray[14][56] ), .D(\bArray[15][56] ), .S0(n8414), .S1(n6993), .Y(
        n6945) );
  CLKINVX1 U14982 ( .A(\xArray[14][57] ), .Y(n8942) );
  CLKINVX1 U14983 ( .A(\xArray[14][58] ), .Y(n8934) );
  CLKINVX1 U14984 ( .A(\xArray[3][59] ), .Y(n8920) );
  CLKINVX1 U14985 ( .A(\xArray[3][60] ), .Y(n8912) );
  MX4X1 U14986 ( .A(\bArray[4][59] ), .B(\bArray[5][59] ), .C(\bArray[6][59] ), 
        .D(\bArray[7][59] ), .S0(n6986), .S1(n6994), .Y(n6959) );
  MX4X1 U14987 ( .A(\bArray[4][58] ), .B(\bArray[5][58] ), .C(\bArray[6][58] ), 
        .D(\bArray[7][58] ), .S0(n6990), .S1(n6994), .Y(n6955) );
  MX4X1 U14988 ( .A(\bArray[4][57] ), .B(\bArray[5][57] ), .C(\bArray[6][57] ), 
        .D(\bArray[7][57] ), .S0(n6990), .S1(n6994), .Y(n6951) );
  MX4X1 U14989 ( .A(\bArray[4][56] ), .B(\bArray[5][56] ), .C(\bArray[6][56] ), 
        .D(\bArray[7][56] ), .S0(n8414), .S1(n6993), .Y(n6947) );
  MX4X1 U14990 ( .A(\bArray[0][56] ), .B(\bArray[1][56] ), .C(\bArray[2][56] ), 
        .D(\bArray[3][56] ), .S0(n7207), .S1(n7212), .Y(n7171) );
  AOI221XL U14991 ( .A0(\xArray[13][56] ), .A1(n8179), .B0(\xArray[1][56] ), 
        .B1(n1747), .C0(n1813), .Y(n1812) );
  OAI22XL U14992 ( .A0(n8175), .A1(n8948), .B0(n8172), .B1(n8946), .Y(n1813)
         );
  AOI221XL U14993 ( .A0(\xArray[13][57] ), .A1(n8179), .B0(\xArray[1][57] ), 
        .B1(n8176), .C0(n1804), .Y(n1803) );
  OAI22XL U14994 ( .A0(n8175), .A1(n8940), .B0(n8172), .B1(n8938), .Y(n1804)
         );
  MX4X1 U14995 ( .A(\bArray[8][57] ), .B(\bArray[9][57] ), .C(\bArray[10][57] ), .D(\bArray[11][57] ), .S0(n7202), .S1(n7213), .Y(n7173) );
  MX4X1 U14996 ( .A(\bArray[12][57] ), .B(\bArray[13][57] ), .C(
        \bArray[14][57] ), .D(\bArray[15][57] ), .S0(n7210), .S1(n7213), .Y(
        n7172) );
  MX4X1 U14997 ( .A(\bArray[4][57] ), .B(\bArray[5][57] ), .C(\bArray[6][57] ), 
        .D(\bArray[7][57] ), .S0(n7202), .S1(n7214), .Y(n7174) );
  MX4X1 U14998 ( .A(\bArray[8][58] ), .B(\bArray[9][58] ), .C(\bArray[10][58] ), .D(\bArray[11][58] ), .S0(n7208), .S1(n7217), .Y(n7177) );
  MX4X1 U14999 ( .A(\bArray[12][58] ), .B(\bArray[13][58] ), .C(
        \bArray[14][58] ), .D(\bArray[15][58] ), .S0(n7211), .S1(n7212), .Y(
        n7176) );
  MX4X1 U15000 ( .A(\bArray[4][58] ), .B(\bArray[5][58] ), .C(\bArray[6][58] ), 
        .D(\bArray[7][58] ), .S0(n7208), .S1(n7222), .Y(n7178) );
  MX4X1 U15001 ( .A(\bArray[8][59] ), .B(\bArray[9][59] ), .C(\bArray[10][59] ), .D(\bArray[11][59] ), .S0(n7201), .S1(N1762), .Y(n7181) );
  MX4X1 U15002 ( .A(\bArray[12][59] ), .B(\bArray[13][59] ), .C(
        \bArray[14][59] ), .D(\bArray[15][59] ), .S0(n7201), .S1(N1762), .Y(
        n7180) );
  MX4X1 U15003 ( .A(\bArray[4][59] ), .B(\bArray[5][59] ), .C(\bArray[6][59] ), 
        .D(\bArray[7][59] ), .S0(n7201), .S1(N1762), .Y(n7182) );
  OAI221X1 U15004 ( .A0(\xArray[7][62] ), .A1(n8289), .B0(\xArray[11][62] ), 
        .B1(n8235), .C0(n984), .Y(n277) );
  OAI221X1 U15005 ( .A0(\xArray[4][62] ), .A1(n8280), .B0(\xArray[8][62] ), 
        .B1(n8226), .C0(n1765), .Y(n1300) );
  OAI221X1 U15006 ( .A0(\xArray[8][62] ), .A1(n8289), .B0(\xArray[12][62] ), 
        .B1(n8235), .C0(n983), .Y(n279) );
  OAI221X1 U15007 ( .A0(\xArray[3][62] ), .A1(n8280), .B0(\xArray[7][62] ), 
        .B1(n8226), .C0(n1764), .Y(n1302) );
  OAI221X1 U15008 ( .A0(\xArray[6][62] ), .A1(n8279), .B0(\xArray[10][62] ), 
        .B1(n8242), .C0(n1303), .Y(n788) );
  OAI221X1 U15009 ( .A0(\xArray[5][62] ), .A1(n8283), .B0(\xArray[9][62] ), 
        .B1(n8229), .C0(n1557), .Y(n982) );
  OA22X1 U15010 ( .A0(\xArray[1][62] ), .A1(n8198), .B0(\xArray[13][62] ), 
        .B1(n8267), .Y(n1557) );
  OAI221XL U15011 ( .A0(\xArray[9][60] ), .A1(n8292), .B0(\xArray[13][60] ), 
        .B1(n8238), .C0(n795), .Y(n294) );
  OA22X1 U15012 ( .A0(\xArray[5][60] ), .A1(n8198), .B0(\xArray[1][60] ), .B1(
        n8254), .Y(n795) );
  OAI221XL U15013 ( .A0(\xArray[2][60] ), .A1(n8280), .B0(\xArray[6][60] ), 
        .B1(n8226), .C0(n1780), .Y(n1562) );
  AOI2BB2X1 U15014 ( .B0(n8918), .B1(n8209), .A0N(\xArray[10][60] ), .A1N(
        n8253), .Y(n1780) );
  OAI222XL U15015 ( .A0(n349), .A1(n8337), .B0(n350), .B1(n8307), .C0(n351), 
        .C1(n7714), .Y(n344) );
  AOI221XL U15016 ( .A0(\xArray[14][53] ), .A1(n6573), .B0(\xArray[2][53] ), 
        .B1(n6579), .C0(n346), .Y(n345) );
  OAI22XL U15017 ( .A0(n8356), .A1(n8971), .B0(n8353), .B1(n8973), .Y(n346) );
  OAI222XL U15018 ( .A0(n357), .A1(n8337), .B0(n358), .B1(n8306), .C0(n359), 
        .C1(n7713), .Y(n352) );
  AOI221XL U15019 ( .A0(\xArray[14][52] ), .A1(n6573), .B0(\xArray[2][52] ), 
        .B1(n8360), .C0(n354), .Y(n353) );
  OAI22XL U15020 ( .A0(n8356), .A1(n8979), .B0(n8353), .B1(n8981), .Y(n354) );
  CLKINVX1 U15021 ( .A(\xArray[14][60] ), .Y(n8918) );
  CLKINVX1 U15022 ( .A(\xArray[14][59] ), .Y(n8926) );
  CLKINVX1 U15023 ( .A(\xArray[5][52] ), .Y(n8978) );
  CLKINVX1 U15024 ( .A(\xArray[5][53] ), .Y(n8970) );
  CLKINVX1 U15025 ( .A(\xArray[5][54] ), .Y(n8962) );
  CLKINVX1 U15026 ( .A(\xArray[5][55] ), .Y(n8954) );
  CLKINVX1 U15027 ( .A(\xArray[3][61] ), .Y(n8904) );
  MX4X1 U15028 ( .A(\bArray[0][57] ), .B(\bArray[1][57] ), .C(\bArray[2][57] ), 
        .D(\bArray[3][57] ), .S0(n7209), .S1(n7215), .Y(n7175) );
  MX4X1 U15029 ( .A(\bArray[0][58] ), .B(\bArray[1][58] ), .C(\bArray[2][58] ), 
        .D(\bArray[3][58] ), .S0(n7201), .S1(N1762), .Y(n7179) );
  MX4X1 U15030 ( .A(\bArray[0][59] ), .B(\bArray[1][59] ), .C(\bArray[2][59] ), 
        .D(\bArray[3][59] ), .S0(n7201), .S1(N1762), .Y(n7183) );
  CLKINVX1 U15031 ( .A(\xArray[9][52] ), .Y(n8980) );
  CLKINVX1 U15032 ( .A(\xArray[9][53] ), .Y(n8972) );
  CLKINVX1 U15033 ( .A(\xArray[9][54] ), .Y(n8964) );
  CLKINVX1 U15034 ( .A(\xArray[9][55] ), .Y(n8956) );
  CLKINVX1 U15035 ( .A(\xArray[6][51] ), .Y(n8987) );
  CLKINVX1 U15036 ( .A(\xArray[6][50] ), .Y(n8995) );
  CLKINVX1 U15037 ( .A(\xArray[6][49] ), .Y(n9003) );
  CLKINVX1 U15038 ( .A(\xArray[6][48] ), .Y(n9011) );
  CLKINVX1 U15039 ( .A(\xArray[10][51] ), .Y(n8989) );
  CLKINVX1 U15040 ( .A(\xArray[10][50] ), .Y(n8997) );
  CLKINVX1 U15041 ( .A(\xArray[10][49] ), .Y(n9005) );
  CLKINVX1 U15042 ( .A(\xArray[10][48] ), .Y(n9013) );
  AOI221XL U15043 ( .A0(\xArray[13][58] ), .A1(n8179), .B0(\xArray[1][58] ), 
        .B1(n8176), .C0(n1795), .Y(n1794) );
  OAI22XL U15044 ( .A0(n8175), .A1(n8932), .B0(n8172), .B1(n8930), .Y(n1795)
         );
  AOI221XL U15045 ( .A0(\xArray[13][59] ), .A1(n8179), .B0(\xArray[1][59] ), 
        .B1(n8176), .C0(n1786), .Y(n1785) );
  OAI22XL U15046 ( .A0(n8175), .A1(n8924), .B0(n8172), .B1(n8922), .Y(n1786)
         );
  MX4X1 U15047 ( .A(\bArray[0][60] ), .B(\bArray[1][60] ), .C(\bArray[2][60] ), 
        .D(\bArray[3][60] ), .S0(n7210), .S1(n7222), .Y(n7187) );
  MX4X1 U15048 ( .A(\bArray[8][60] ), .B(\bArray[9][60] ), .C(\bArray[10][60] ), .D(\bArray[11][60] ), .S0(n7201), .S1(n7222), .Y(n7185) );
  MX4X1 U15049 ( .A(\bArray[12][60] ), .B(\bArray[13][60] ), .C(
        \bArray[14][60] ), .D(\bArray[15][60] ), .S0(n7201), .S1(n7222), .Y(
        n7184) );
  MX4X1 U15050 ( .A(\bArray[8][61] ), .B(\bArray[9][61] ), .C(\bArray[10][61] ), .D(\bArray[11][61] ), .S0(n7202), .S1(n7214), .Y(n7189) );
  MX4X1 U15051 ( .A(\bArray[12][61] ), .B(\bArray[13][61] ), .C(
        \bArray[14][61] ), .D(\bArray[15][61] ), .S0(n7202), .S1(n7222), .Y(
        n7188) );
  MX4X1 U15052 ( .A(\bArray[4][61] ), .B(\bArray[5][61] ), .C(\bArray[6][61] ), 
        .D(\bArray[7][61] ), .S0(n7202), .S1(n7214), .Y(n7190) );
  MX4X1 U15053 ( .A(\bArray[8][62] ), .B(\bArray[9][62] ), .C(\bArray[10][62] ), .D(\bArray[11][62] ), .S0(n7210), .S1(n8409), .Y(n7193) );
  MX4X1 U15054 ( .A(\bArray[12][62] ), .B(\bArray[13][62] ), .C(
        \bArray[14][62] ), .D(\bArray[15][62] ), .S0(n7202), .S1(n8409), .Y(
        n7192) );
  MX4X1 U15055 ( .A(\bArray[4][62] ), .B(\bArray[5][62] ), .C(\bArray[6][62] ), 
        .D(\bArray[7][62] ), .S0(n7210), .S1(n8409), .Y(n7194) );
  OAI221XL U15056 ( .A0(\xArray[9][61] ), .A1(n8292), .B0(\xArray[13][61] ), 
        .B1(n8238), .C0(n792), .Y(n286) );
  OA22X1 U15057 ( .A0(\xArray[5][61] ), .A1(n8198), .B0(\xArray[1][61] ), .B1(
        n8258), .Y(n792) );
  OAI221XL U15058 ( .A0(\xArray[9][62] ), .A1(n8292), .B0(\xArray[13][62] ), 
        .B1(n8238), .C0(n789), .Y(n278) );
  OA22X1 U15059 ( .A0(\xArray[5][62] ), .A1(n786), .B0(\xArray[1][62] ), .B1(
        n8254), .Y(n789) );
  OAI221XL U15060 ( .A0(\xArray[2][61] ), .A1(n8280), .B0(\xArray[6][61] ), 
        .B1(n8226), .C0(n1771), .Y(n1559) );
  AOI2BB2X1 U15061 ( .B0(n8910), .B1(n8209), .A0N(\xArray[10][61] ), .A1N(
        n8253), .Y(n1771) );
  OAI221XL U15062 ( .A0(\xArray[2][62] ), .A1(n8280), .B0(\xArray[6][62] ), 
        .B1(n8226), .C0(n1762), .Y(n1556) );
  OAI222XL U15063 ( .A0(n333), .A1(n8337), .B0(n334), .B1(n8310), .C0(n335), 
        .C1(n7714), .Y(n328) );
  AOI221XL U15064 ( .A0(\xArray[14][55] ), .A1(n6573), .B0(\xArray[2][55] ), 
        .B1(n6579), .C0(n330), .Y(n329) );
  OAI22XL U15065 ( .A0(n8359), .A1(n8955), .B0(n8353), .B1(n8957), .Y(n330) );
  OAI222XL U15066 ( .A0(n341), .A1(n8337), .B0(n342), .B1(n8320), .C0(n343), 
        .C1(n7714), .Y(n336) );
  AOI221XL U15067 ( .A0(\xArray[14][54] ), .A1(n6573), .B0(\xArray[2][54] ), 
        .B1(n6579), .C0(n338), .Y(n337) );
  OAI22XL U15068 ( .A0(n8356), .A1(n8963), .B0(n8353), .B1(n8965), .Y(n338) );
  MX4X1 U15069 ( .A(n6968), .B(n6966), .C(n6967), .D(n6965), .S0(n7007), .S1(
        N1759), .Y(N25539) );
  MX4X1 U15070 ( .A(\bArray[8][61] ), .B(\bArray[9][61] ), .C(\bArray[10][61] ), .D(\bArray[11][61] ), .S0(n6978), .S1(n7001), .Y(n6966) );
  MX4X1 U15071 ( .A(\bArray[0][61] ), .B(\bArray[1][61] ), .C(\bArray[2][61] ), 
        .D(\bArray[3][61] ), .S0(n6978), .S1(n7000), .Y(n6968) );
  MX4X1 U15072 ( .A(\bArray[12][61] ), .B(\bArray[13][61] ), .C(
        \bArray[14][61] ), .D(\bArray[15][61] ), .S0(n6978), .S1(n6991), .Y(
        n6965) );
  MX4X1 U15073 ( .A(n6964), .B(n6962), .C(n6963), .D(n6961), .S0(n7007), .S1(
        N1759), .Y(N25540) );
  MX4X1 U15074 ( .A(\bArray[0][60] ), .B(\bArray[1][60] ), .C(\bArray[2][60] ), 
        .D(\bArray[3][60] ), .S0(n6978), .S1(n6993), .Y(n6964) );
  MX4X1 U15075 ( .A(\bArray[8][60] ), .B(\bArray[9][60] ), .C(\bArray[10][60] ), .D(\bArray[11][60] ), .S0(n6977), .S1(n6993), .Y(n6962) );
  MX4X1 U15076 ( .A(\bArray[12][60] ), .B(\bArray[13][60] ), .C(
        \bArray[14][60] ), .D(\bArray[15][60] ), .S0(n6985), .S1(n6993), .Y(
        n6961) );
  MX4X1 U15077 ( .A(n6972), .B(n6970), .C(n6971), .D(n6969), .S0(n7007), .S1(
        N1759), .Y(N25538) );
  MX4X1 U15078 ( .A(\bArray[8][62] ), .B(\bArray[9][62] ), .C(\bArray[10][62] ), .D(\bArray[11][62] ), .S0(n6979), .S1(n6995), .Y(n6970) );
  MX4X1 U15079 ( .A(\bArray[0][62] ), .B(\bArray[1][62] ), .C(\bArray[2][62] ), 
        .D(\bArray[3][62] ), .S0(n6979), .S1(n6995), .Y(n6972) );
  MX4X1 U15080 ( .A(\bArray[12][62] ), .B(\bArray[13][62] ), .C(
        \bArray[14][62] ), .D(\bArray[15][62] ), .S0(n6979), .S1(n6994), .Y(
        n6969) );
  MX4X1 U15081 ( .A(n6976), .B(n6974), .C(n6975), .D(n6973), .S0(n7007), .S1(
        n8412), .Y(n6784) );
  MX4X1 U15082 ( .A(\bArray[8][63] ), .B(\bArray[9][63] ), .C(\bArray[10][63] ), .D(\bArray[11][63] ), .S0(n6978), .S1(n6992), .Y(n6974) );
  MX4X1 U15083 ( .A(\bArray[0][63] ), .B(\bArray[1][63] ), .C(\bArray[2][63] ), 
        .D(\bArray[3][63] ), .S0(n6978), .S1(n6992), .Y(n6976) );
  MX4X1 U15084 ( .A(\bArray[12][63] ), .B(\bArray[13][63] ), .C(
        \bArray[14][63] ), .D(\bArray[15][63] ), .S0(n6978), .S1(n7001), .Y(
        n6973) );
  CLKINVX1 U15085 ( .A(\xArray[14][61] ), .Y(n8910) );
  CLKINVX1 U15086 ( .A(\xArray[3][62] ), .Y(n8896) );
  MX4X1 U15087 ( .A(\bArray[4][61] ), .B(\bArray[5][61] ), .C(\bArray[6][61] ), 
        .D(\bArray[7][61] ), .S0(n6978), .S1(n7002), .Y(n6967) );
  MX4X1 U15088 ( .A(\bArray[4][60] ), .B(\bArray[5][60] ), .C(\bArray[6][60] ), 
        .D(\bArray[7][60] ), .S0(n6978), .S1(n6993), .Y(n6963) );
  MX4X1 U15089 ( .A(\bArray[4][62] ), .B(\bArray[5][62] ), .C(\bArray[6][62] ), 
        .D(\bArray[7][62] ), .S0(n6978), .S1(n6999), .Y(n6971) );
  MX4X1 U15090 ( .A(\bArray[4][60] ), .B(\bArray[5][60] ), .C(\bArray[6][60] ), 
        .D(\bArray[7][60] ), .S0(n7203), .S1(n7222), .Y(n7186) );
  MX4X1 U15091 ( .A(\bArray[4][63] ), .B(\bArray[5][63] ), .C(\bArray[6][63] ), 
        .D(\bArray[7][63] ), .S0(n6986), .S1(n6993), .Y(n6975) );
  MX4X1 U15092 ( .A(\bArray[0][61] ), .B(\bArray[1][61] ), .C(\bArray[2][61] ), 
        .D(\bArray[3][61] ), .S0(n7202), .S1(n7222), .Y(n7191) );
  MX4X1 U15093 ( .A(\bArray[0][62] ), .B(\bArray[1][62] ), .C(\bArray[2][62] ), 
        .D(\bArray[3][62] ), .S0(n7202), .S1(N1762), .Y(n7195) );
  CLKINVX1 U15094 ( .A(\xArray[10][52] ), .Y(n8981) );
  AOI221XL U15095 ( .A0(\xArray[13][60] ), .A1(n8179), .B0(\xArray[1][60] ), 
        .B1(n8176), .C0(n1777), .Y(n1776) );
  OAI22XL U15096 ( .A0(n8175), .A1(n8916), .B0(n8170), .B1(n8914), .Y(n1777)
         );
  AOI221XL U15097 ( .A0(\xArray[13][61] ), .A1(n8181), .B0(\xArray[1][61] ), 
        .B1(n8176), .C0(n1768), .Y(n1767) );
  OAI22XL U15098 ( .A0(n8175), .A1(n8908), .B0(n8170), .B1(n8906), .Y(n1768)
         );
  AOI221XL U15099 ( .A0(\xArray[13][62] ), .A1(n8180), .B0(\xArray[1][62] ), 
        .B1(n8176), .C0(n1759), .Y(n1758) );
  OAI22XL U15100 ( .A0(n8175), .A1(n8900), .B0(n8170), .B1(n8898), .Y(n1759)
         );
  MX4X1 U15101 ( .A(\bArray[8][63] ), .B(\bArray[9][63] ), .C(\bArray[10][63] ), .D(\bArray[11][63] ), .S0(n7204), .S1(n8409), .Y(n7197) );
  MX4X1 U15102 ( .A(\bArray[12][63] ), .B(\bArray[13][63] ), .C(
        \bArray[14][63] ), .D(\bArray[15][63] ), .S0(n7204), .S1(n8409), .Y(
        n7196) );
  MX4X1 U15103 ( .A(\bArray[4][63] ), .B(\bArray[5][63] ), .C(\bArray[6][63] ), 
        .D(\bArray[7][63] ), .S0(n7202), .S1(n8409), .Y(n7198) );
  OAI221X1 U15104 ( .A0(\xArray[7][63] ), .A1(n8289), .B0(\xArray[11][63] ), 
        .B1(n8235), .C0(n979), .Y(n267) );
  OAI221X1 U15105 ( .A0(\xArray[4][63] ), .A1(n8280), .B0(\xArray[8][63] ), 
        .B1(n8226), .C0(n1756), .Y(n1296) );
  OAI221X1 U15106 ( .A0(\xArray[8][63] ), .A1(n8289), .B0(\xArray[12][63] ), 
        .B1(n8235), .C0(n978), .Y(n271) );
  OAI221X1 U15107 ( .A0(\xArray[6][63] ), .A1(n8295), .B0(\xArray[10][63] ), 
        .B1(n8241), .C0(n1299), .Y(n784) );
  OAI221X1 U15108 ( .A0(\xArray[3][63] ), .A1(n8280), .B0(\xArray[7][63] ), 
        .B1(n8226), .C0(n1755), .Y(n1298) );
  OAI221X1 U15109 ( .A0(\xArray[5][63] ), .A1(n8279), .B0(\xArray[9][63] ), 
        .B1(n8242), .C0(n1554), .Y(n977) );
  OAI222XL U15110 ( .A0(n309), .A1(n8337), .B0(n310), .B1(n8309), .C0(n311), 
        .C1(n7714), .Y(n304) );
  AOI221XL U15111 ( .A0(\xArray[14][58] ), .A1(n6573), .B0(\xArray[2][58] ), 
        .B1(n8362), .C0(n306), .Y(n305) );
  OAI22XL U15112 ( .A0(n8359), .A1(n8931), .B0(n8353), .B1(n8933), .Y(n306) );
  OAI222XL U15113 ( .A0(n317), .A1(n8337), .B0(n318), .B1(n8311), .C0(n319), 
        .C1(n7714), .Y(n312) );
  AOI221XL U15114 ( .A0(\xArray[14][57] ), .A1(n6573), .B0(\xArray[2][57] ), 
        .B1(n6579), .C0(n314), .Y(n313) );
  OAI22XL U15115 ( .A0(n8359), .A1(n8939), .B0(n8353), .B1(n8941), .Y(n314) );
  OAI222XL U15116 ( .A0(n325), .A1(n8337), .B0(n326), .B1(n8310), .C0(n327), 
        .C1(n7714), .Y(n320) );
  AOI221XL U15117 ( .A0(\xArray[14][56] ), .A1(n6573), .B0(\xArray[2][56] ), 
        .B1(n6579), .C0(n322), .Y(n321) );
  OAI22XL U15118 ( .A0(n8359), .A1(n8947), .B0(n8353), .B1(n8949), .Y(n322) );
  CLKINVX1 U15119 ( .A(\xArray[14][62] ), .Y(n8902) );
  CLKINVX1 U15120 ( .A(\xArray[5][56] ), .Y(n8946) );
  CLKINVX1 U15121 ( .A(\xArray[5][57] ), .Y(n8938) );
  CLKINVX1 U15122 ( .A(\xArray[5][58] ), .Y(n8930) );
  CLKINVX1 U15123 ( .A(\xArray[5][59] ), .Y(n8922) );
  MX4X1 U15124 ( .A(\bArray[0][63] ), .B(\bArray[1][63] ), .C(\bArray[2][63] ), 
        .D(\bArray[3][63] ), .S0(N1761), .S1(n8409), .Y(n7199) );
  CLKINVX1 U15125 ( .A(\xArray[9][56] ), .Y(n8948) );
  CLKINVX1 U15126 ( .A(\xArray[9][57] ), .Y(n8940) );
  CLKINVX1 U15127 ( .A(\xArray[9][58] ), .Y(n8932) );
  CLKINVX1 U15128 ( .A(\xArray[9][59] ), .Y(n8924) );
  CLKINVX1 U15129 ( .A(\xArray[6][55] ), .Y(n8955) );
  CLKINVX1 U15130 ( .A(\xArray[6][54] ), .Y(n8963) );
  CLKINVX1 U15131 ( .A(\xArray[6][53] ), .Y(n8971) );
  CLKINVX1 U15132 ( .A(\xArray[6][52] ), .Y(n8979) );
  CLKINVX1 U15133 ( .A(\xArray[10][55] ), .Y(n8957) );
  CLKINVX1 U15134 ( .A(\xArray[10][54] ), .Y(n8965) );
  CLKINVX1 U15135 ( .A(\xArray[10][53] ), .Y(n8973) );
  AOI221XL U15136 ( .A0(\xArray[13][63] ), .A1(n8181), .B0(\xArray[1][63] ), 
        .B1(n8176), .C0(n1748), .Y(n1745) );
  OAI22XL U15137 ( .A0(n1749), .A1(n8892), .B0(n8170), .B1(n8890), .Y(n1748)
         );
  OAI221XL U15138 ( .A0(\xArray[2][63] ), .A1(n8280), .B0(\xArray[6][63] ), 
        .B1(n8226), .C0(n1753), .Y(n1553) );
  OAI222XL U15139 ( .A0(n301), .A1(n8337), .B0(n302), .B1(n8318), .C0(n303), 
        .C1(n7717), .Y(n296) );
  AOI221XL U15140 ( .A0(\xArray[14][59] ), .A1(n6573), .B0(\xArray[2][59] ), 
        .B1(n8362), .C0(n298), .Y(n297) );
  OAI22XL U15141 ( .A0(n8359), .A1(n8923), .B0(n8353), .B1(n8925), .Y(n298) );
  CLKINVX1 U15142 ( .A(\xArray[5][60] ), .Y(n8914) );
  CLKINVX1 U15143 ( .A(\xArray[5][61] ), .Y(n8906) );
  CLKINVX1 U15144 ( .A(\xArray[3][63] ), .Y(n8888) );
  CLKINVX1 U15145 ( .A(\xArray[9][60] ), .Y(n8916) );
  CLKINVX1 U15146 ( .A(\xArray[9][61] ), .Y(n8908) );
  CLKINVX1 U15147 ( .A(\xArray[6][56] ), .Y(n8947) );
  CLKINVX1 U15148 ( .A(\xArray[10][56] ), .Y(n8949) );
  OAI221XL U15149 ( .A0(\xArray[9][63] ), .A1(n8279), .B0(\xArray[13][63] ), 
        .B1(n8225), .C0(n785), .Y(n269) );
  OAI222XL U15150 ( .A0(n293), .A1(n8337), .B0(n294), .B1(n8309), .C0(n295), 
        .C1(n7729), .Y(n288) );
  AOI221XL U15151 ( .A0(\xArray[14][60] ), .A1(n6573), .B0(\xArray[2][60] ), 
        .B1(n8362), .C0(n290), .Y(n289) );
  OAI22XL U15152 ( .A0(n8356), .A1(n8915), .B0(n8353), .B1(n8917), .Y(n290) );
  OAI222XL U15153 ( .A0(n285), .A1(n8337), .B0(n286), .B1(n8309), .C0(n287), 
        .C1(n7720), .Y(n280) );
  AOI221XL U15154 ( .A0(\xArray[14][61] ), .A1(n6573), .B0(\xArray[2][61] ), 
        .B1(n8362), .C0(n282), .Y(n281) );
  OAI22XL U15155 ( .A0(n8356), .A1(n8907), .B0(n8353), .B1(n8909), .Y(n282) );
  OAI222XL U15156 ( .A0(n277), .A1(n8337), .B0(n278), .B1(n8309), .C0(n279), 
        .C1(n7729), .Y(n272) );
  AOI221XL U15157 ( .A0(\xArray[14][62] ), .A1(n6573), .B0(\xArray[2][62] ), 
        .B1(n8362), .C0(n274), .Y(n273) );
  OAI22XL U15158 ( .A0(n8356), .A1(n8899), .B0(n8353), .B1(n8901), .Y(n274) );
  OAI222XL U15159 ( .A0(n8340), .A1(n267), .B0(n8320), .B1(n269), .C0(n7713), 
        .C1(n271), .Y(n257) );
  AOI221XL U15160 ( .A0(\xArray[14][63] ), .A1(n6573), .B0(\xArray[2][63] ), 
        .B1(n8362), .C0(n261), .Y(n258) );
  OAI22XL U15161 ( .A0(n8356), .A1(n8891), .B0(n8353), .B1(n8893), .Y(n261) );
  CLKINVX1 U15162 ( .A(\xArray[14][63] ), .Y(n8894) );
  CLKINVX1 U15163 ( .A(\xArray[5][62] ), .Y(n8898) );
  CLKINVX1 U15164 ( .A(\xArray[5][63] ), .Y(n8890) );
  CLKINVX1 U15165 ( .A(\xArray[9][62] ), .Y(n8900) );
  CLKINVX1 U15166 ( .A(\xArray[9][63] ), .Y(n8892) );
  CLKINVX1 U15167 ( .A(\xArray[6][59] ), .Y(n8923) );
  CLKINVX1 U15168 ( .A(\xArray[6][58] ), .Y(n8931) );
  CLKINVX1 U15169 ( .A(\xArray[6][57] ), .Y(n8939) );
  CLKINVX1 U15170 ( .A(\xArray[10][59] ), .Y(n8925) );
  CLKINVX1 U15171 ( .A(\xArray[10][58] ), .Y(n8933) );
  CLKINVX1 U15172 ( .A(\xArray[10][57] ), .Y(n8941) );
  CLKINVX1 U15173 ( .A(\xArray[6][60] ), .Y(n8915) );
  CLKINVX1 U15174 ( .A(\xArray[6][61] ), .Y(n8907) );
  CLKINVX1 U15175 ( .A(\xArray[6][62] ), .Y(n8899) );
  CLKINVX1 U15176 ( .A(\xArray[10][60] ), .Y(n8917) );
  CLKINVX1 U15177 ( .A(\xArray[10][61] ), .Y(n8909) );
  CLKINVX1 U15178 ( .A(\xArray[10][62] ), .Y(n8901) );
  CLKINVX1 U15179 ( .A(\xArray[6][63] ), .Y(n8891) );
  CLKINVX1 U15180 ( .A(\xArray[10][63] ), .Y(n8893) );
  AND2X2 U15181 ( .A(N1804), .B(n8405), .Y(N1837) );
  NOR2X1 U15182 ( .A(n6736), .B(n102), .Y(n4831) );
  OR2X1 U15183 ( .A(n8425), .B(n8424), .Y(n6736) );
  NOR4X1 U15184 ( .A(n4879), .B(xCount[31]), .C(xCount[5]), .D(xCount[4]), .Y(
        n4878) );
  NAND4X1 U15185 ( .A(n109), .B(n110), .C(n111), .D(n112), .Y(n4879) );
  AND4X1 U15186 ( .A(n4875), .B(n4876), .C(n4877), .D(n4878), .Y(n4867) );
  NOR4X1 U15187 ( .A(n4882), .B(xCount[10]), .C(xCount[12]), .D(xCount[11]), 
        .Y(n4875) );
  NOR4X1 U15188 ( .A(n4881), .B(xCount[17]), .C(xCount[19]), .D(xCount[18]), 
        .Y(n4876) );
  NOR4X1 U15189 ( .A(n4880), .B(xCount[24]), .C(xCount[26]), .D(xCount[25]), 
        .Y(n4877) );
  OAI2BB2XL U15190 ( .B0(n4902), .B1(n8400), .A0N(N35048), .A1N(n8395), .Y(
        n5707) );
  OAI2BB2XL U15191 ( .B0(n4903), .B1(n8400), .A0N(N35047), .A1N(n8395), .Y(
        n5708) );
  OAI2BB2XL U15192 ( .B0(n4904), .B1(n8400), .A0N(N35046), .A1N(n8395), .Y(
        n5709) );
  OAI2BB2XL U15193 ( .B0(n4905), .B1(n8400), .A0N(N35045), .A1N(n8395), .Y(
        n5710) );
  OAI2BB2XL U15194 ( .B0(n4906), .B1(n8400), .A0N(N35044), .A1N(n8395), .Y(
        n5711) );
  NOR2BX1 U15195 ( .AN(N35115), .B(n8398), .Y(outCount_next[31]) );
  NAND4X1 U15196 ( .A(n130), .B(n131), .C(n132), .D(n133), .Y(n4880) );
  NAND4X1 U15197 ( .A(n123), .B(n124), .C(n125), .D(n126), .Y(n4881) );
  NAND4X1 U15198 ( .A(n116), .B(n117), .C(n118), .D(n119), .Y(n4882) );
  OAI2BB2XL U15199 ( .B0(n4907), .B1(n8400), .A0N(N35043), .A1N(n8396), .Y(
        n5712) );
  OAI2BB2XL U15200 ( .B0(n4908), .B1(n8400), .A0N(N35042), .A1N(n8396), .Y(
        n5713) );
  OAI2BB2XL U15201 ( .B0(n4909), .B1(n8399), .A0N(N35041), .A1N(n8396), .Y(
        n5714) );
  OAI2BB2XL U15202 ( .B0(n4910), .B1(n8400), .A0N(N35040), .A1N(n8396), .Y(
        n5715) );
  OAI2BB2XL U15203 ( .B0(n4911), .B1(n8399), .A0N(N35039), .A1N(n8396), .Y(
        n5716) );
  OAI2BB2XL U15204 ( .B0(n4912), .B1(n8399), .A0N(N35038), .A1N(n8396), .Y(
        n5717) );
  OAI2BB2XL U15205 ( .B0(n4913), .B1(n8399), .A0N(N35037), .A1N(n8396), .Y(
        n5718) );
  OAI211X1 U15206 ( .A0(n102), .A1(n241), .B0(n8398), .C0(n161), .Y(
        state_next[1]) );
  OAI211X1 U15207 ( .A0(n242), .A1(n243), .B0(n8398), .C0(n244), .Y(
        state_next[0]) );
  NAND4X1 U15208 ( .A(n248), .B(n249), .C(n250), .D(n251), .Y(n243) );
  NAND4BX1 U15209 ( .AN(n252), .B(n253), .C(n254), .D(n255), .Y(n242) );
  AOI32X1 U15210 ( .A0(n6624), .A1(n6620), .A2(n8405), .B0(n102), .B1(n8854), 
        .Y(n244) );
  NAND3BX1 U15211 ( .AN(n6737), .B(state[1]), .C(state[0]), .Y(n159) );
  OR2X1 U15212 ( .A(n8447), .B(n8446), .Y(n6737) );
  NOR4X1 U15213 ( .A(n4884), .B(n4885), .C(n4886), .D(n4887), .Y(n3148) );
  NAND4BX1 U15214 ( .AN(n4891), .B(n101), .C(n99), .D(n100), .Y(n4884) );
  NAND4BX1 U15215 ( .AN(n4890), .B(n94), .C(n92), .D(n93), .Y(n4885) );
  NAND4BX1 U15216 ( .AN(n4889), .B(n87), .C(n85), .D(n86), .Y(n4886) );
  NAND4BX1 U15217 ( .AN(n4888), .B(n80), .C(n78), .D(n79), .Y(n4887) );
  NAND4X1 U15218 ( .A(n77), .B(n76), .C(n75), .D(n73), .Y(n4888) );
  NOR2BX1 U15219 ( .AN(n3148), .B(n74), .Y(n3638) );
  OAI2BB2XL U15220 ( .B0(n4920), .B1(n8399), .A0N(N35030), .A1N(n8395), .Y(
        n5725) );
  OAI2BB2XL U15221 ( .B0(n4923), .B1(n8399), .A0N(N35027), .A1N(n8396), .Y(
        n5728) );
  OAI2BB2XL U15222 ( .B0(n4914), .B1(n8399), .A0N(N35036), .A1N(n8396), .Y(
        n5719) );
  OAI2BB2XL U15223 ( .B0(n4915), .B1(n8399), .A0N(N35035), .A1N(n8396), .Y(
        n5720) );
  OAI2BB2XL U15224 ( .B0(n4916), .B1(n8399), .A0N(N35034), .A1N(n8396), .Y(
        n5721) );
  OAI2BB2XL U15225 ( .B0(n4917), .B1(n8399), .A0N(N35033), .A1N(n8396), .Y(
        n5722) );
  OAI2BB2XL U15226 ( .B0(n4918), .B1(n8399), .A0N(N35032), .A1N(n8396), .Y(
        n5723) );
  OAI2BB2XL U15227 ( .B0(n4919), .B1(n8399), .A0N(N35031), .A1N(n160), .Y(
        n5724) );
  OAI2BB2XL U15228 ( .B0(n4921), .B1(n8399), .A0N(N35029), .A1N(n160), .Y(
        n5726) );
  OAI2BB2XL U15229 ( .B0(n4922), .B1(n8399), .A0N(N35028), .A1N(n160), .Y(
        n5727) );
  OAI2BB2XL U15230 ( .B0(n4926), .B1(n8400), .A0N(N35024), .A1N(n8395), .Y(
        n5731) );
  OAI2BB2XL U15231 ( .B0(n4927), .B1(n8400), .A0N(N35023), .A1N(n8395), .Y(
        n5732) );
  OAI2BB2XL U15232 ( .B0(n4928), .B1(n8400), .A0N(N35022), .A1N(n8395), .Y(
        n5733) );
  OAI2BB2XL U15233 ( .B0(n4929), .B1(n8400), .A0N(N35021), .A1N(n8395), .Y(
        n5734) );
  OAI2BB2XL U15234 ( .B0(n4930), .B1(n8400), .A0N(N35020), .A1N(n8395), .Y(
        n5735) );
  OAI2BB2XL U15235 ( .B0(n4931), .B1(n8400), .A0N(N35019), .A1N(n8395), .Y(
        n5736) );
  OAI2BB2XL U15236 ( .B0(n4932), .B1(n8401), .A0N(N35018), .A1N(n8396), .Y(
        n5737) );
  OAI2BB2XL U15237 ( .B0(n4933), .B1(n8401), .A0N(N35017), .A1N(n160), .Y(
        n5738) );
  OAI2BB2XL U15238 ( .B0(n4924), .B1(n8401), .A0N(N35026), .A1N(n8395), .Y(
        n5729) );
  OAI2BB2XL U15239 ( .B0(n4925), .B1(n8401), .A0N(N35025), .A1N(n8395), .Y(
        n5730) );
  AND2X2 U15240 ( .A(N34941), .B(n8403), .Y(N34942) );
  MX4X1 U15241 ( .A(n7231), .B(n7229), .C(n7230), .D(n7228), .S0(n7356), .S1(
        n7359), .Y(N34941) );
  AND2X2 U15242 ( .A(N34940), .B(n8402), .Y(N34943) );
  MX4X1 U15243 ( .A(n7235), .B(n7233), .C(n7234), .D(n7232), .S0(n7356), .S1(
        n7360), .Y(N34940) );
  OAI21XL U15244 ( .A0(n4972), .A1(n7699), .B0(n8375), .Y(n5777) );
  OAI21XL U15245 ( .A0(n4973), .A1(n7699), .B0(n8375), .Y(n5778) );
  OAI21XL U15246 ( .A0(n4974), .A1(n7699), .B0(n8375), .Y(n5779) );
  OAI21XL U15247 ( .A0(n4975), .A1(n7699), .B0(n8375), .Y(n5780) );
  OAI21XL U15248 ( .A0(n4976), .A1(n7699), .B0(n8375), .Y(n5781) );
  OAI21XL U15249 ( .A0(n4977), .A1(n6719), .B0(n8375), .Y(n5782) );
  OAI21XL U15250 ( .A0(n4978), .A1(n6719), .B0(n8375), .Y(n5783) );
  OAI21XL U15251 ( .A0(n4979), .A1(n6719), .B0(n8375), .Y(n5784) );
  OAI21XL U15252 ( .A0(n4980), .A1(n6719), .B0(n8375), .Y(n5785) );
  OAI21XL U15253 ( .A0(n5020), .A1(n7686), .B0(n8373), .Y(n5825) );
  OAI21XL U15254 ( .A0(n5021), .A1(n7686), .B0(n8373), .Y(n5826) );
  OAI21XL U15255 ( .A0(n5022), .A1(n7686), .B0(n8373), .Y(n5827) );
  OAI21XL U15256 ( .A0(n5023), .A1(n7686), .B0(n8373), .Y(n5828) );
  OAI21XL U15257 ( .A0(n5024), .A1(n7687), .B0(n8373), .Y(n5829) );
  OAI21XL U15258 ( .A0(n5025), .A1(n7687), .B0(n8373), .Y(n5830) );
  OAI21XL U15259 ( .A0(n5026), .A1(n7687), .B0(n8373), .Y(n5831) );
  OAI21XL U15260 ( .A0(n5027), .A1(n7687), .B0(n8373), .Y(n5832) );
  OAI21XL U15261 ( .A0(n5028), .A1(n7687), .B0(n8373), .Y(n5833) );
  OAI21XL U15262 ( .A0(n5068), .A1(n7689), .B0(n8371), .Y(n5873) );
  OAI21XL U15263 ( .A0(n5069), .A1(n7689), .B0(n8371), .Y(n5874) );
  OAI21XL U15264 ( .A0(n5070), .A1(n7689), .B0(n8371), .Y(n5875) );
  OAI21XL U15265 ( .A0(n5071), .A1(n7689), .B0(n8371), .Y(n5876) );
  OAI21XL U15266 ( .A0(n5072), .A1(n7689), .B0(n8371), .Y(n5877) );
  OAI21XL U15267 ( .A0(n5073), .A1(n6721), .B0(n8371), .Y(n5878) );
  OAI21XL U15268 ( .A0(n5074), .A1(n6721), .B0(n8371), .Y(n5879) );
  OAI21XL U15269 ( .A0(n5075), .A1(n6721), .B0(n8371), .Y(n5880) );
  OAI21XL U15270 ( .A0(n5076), .A1(n6721), .B0(n8371), .Y(n5881) );
  OAI21XL U15271 ( .A0(n5116), .A1(n7690), .B0(n8369), .Y(n5921) );
  OAI21XL U15272 ( .A0(n5117), .A1(n7690), .B0(n8369), .Y(n5922) );
  OAI21XL U15273 ( .A0(n5118), .A1(n7690), .B0(n8369), .Y(n5923) );
  OAI21XL U15274 ( .A0(n5119), .A1(n7691), .B0(n8369), .Y(n5924) );
  OAI21XL U15275 ( .A0(n5120), .A1(n7691), .B0(n8369), .Y(n5925) );
  OAI21XL U15276 ( .A0(n5121), .A1(n7691), .B0(n8369), .Y(n5926) );
  OAI21XL U15277 ( .A0(n5122), .A1(n7691), .B0(n8369), .Y(n5927) );
  OAI21XL U15278 ( .A0(n5123), .A1(n7691), .B0(n8369), .Y(n5928) );
  OAI21XL U15279 ( .A0(n5124), .A1(n7691), .B0(n8369), .Y(n5929) );
  OAI21XL U15280 ( .A0(n5164), .A1(n7693), .B0(n8367), .Y(n5969) );
  OAI21XL U15281 ( .A0(n5165), .A1(n7693), .B0(n8367), .Y(n5970) );
  OAI21XL U15282 ( .A0(n5166), .A1(n7693), .B0(n8367), .Y(n5971) );
  OAI21XL U15283 ( .A0(n5167), .A1(n7693), .B0(n8367), .Y(n5972) );
  OAI21XL U15284 ( .A0(n5168), .A1(n7693), .B0(n8367), .Y(n5973) );
  OAI21XL U15285 ( .A0(n5169), .A1(n6723), .B0(n8367), .Y(n5974) );
  OAI21XL U15286 ( .A0(n5170), .A1(n6723), .B0(n8367), .Y(n5975) );
  OAI21XL U15287 ( .A0(n5171), .A1(n6723), .B0(n8367), .Y(n5976) );
  OAI21XL U15288 ( .A0(n5172), .A1(n6723), .B0(n8367), .Y(n5977) );
  OAI21XL U15289 ( .A0(n5212), .A1(n7695), .B0(n8365), .Y(n6017) );
  OAI21XL U15290 ( .A0(n5213), .A1(n7695), .B0(n8365), .Y(n6018) );
  OAI21XL U15291 ( .A0(n5214), .A1(n7695), .B0(n8365), .Y(n6019) );
  OAI21XL U15292 ( .A0(n5215), .A1(n7695), .B0(n8365), .Y(n6020) );
  OAI21XL U15293 ( .A0(n5216), .A1(n7695), .B0(n8365), .Y(n6021) );
  OAI21XL U15294 ( .A0(n5217), .A1(n6724), .B0(n8365), .Y(n6022) );
  OAI21XL U15295 ( .A0(n5218), .A1(n6724), .B0(n8365), .Y(n6023) );
  OAI21XL U15296 ( .A0(n5219), .A1(n6724), .B0(n8365), .Y(n6024) );
  OAI21XL U15297 ( .A0(n5220), .A1(n6724), .B0(n8365), .Y(n6025) );
  OAI21XL U15298 ( .A0(n5260), .A1(n7669), .B0(n8393), .Y(n6065) );
  OAI21XL U15299 ( .A0(n5261), .A1(n7669), .B0(n8393), .Y(n6066) );
  OAI21XL U15300 ( .A0(n5262), .A1(n7669), .B0(n8393), .Y(n6067) );
  OAI21XL U15301 ( .A0(n5263), .A1(n7669), .B0(n8393), .Y(n6068) );
  OAI21XL U15302 ( .A0(n5264), .A1(n7669), .B0(n8393), .Y(n6069) );
  OAI21XL U15303 ( .A0(n5265), .A1(n6734), .B0(n8393), .Y(n6070) );
  OAI21XL U15304 ( .A0(n5266), .A1(n6734), .B0(n8393), .Y(n6071) );
  OAI21XL U15305 ( .A0(n5267), .A1(n6734), .B0(n8393), .Y(n6072) );
  OAI21XL U15306 ( .A0(n5268), .A1(n6734), .B0(n8393), .Y(n6073) );
  OAI21XL U15307 ( .A0(n5308), .A1(n7671), .B0(n8391), .Y(n6113) );
  OAI21XL U15308 ( .A0(n5309), .A1(n7671), .B0(n8391), .Y(n6114) );
  OAI21XL U15309 ( .A0(n5310), .A1(n7671), .B0(n8391), .Y(n6115) );
  OAI21XL U15310 ( .A0(n5311), .A1(n7671), .B0(n8391), .Y(n6116) );
  OAI21XL U15311 ( .A0(n5312), .A1(n7671), .B0(n8391), .Y(n6117) );
  OAI21XL U15312 ( .A0(n5313), .A1(n6725), .B0(n8391), .Y(n6118) );
  OAI21XL U15313 ( .A0(n5314), .A1(n6725), .B0(n8391), .Y(n6119) );
  OAI21XL U15314 ( .A0(n5315), .A1(n6725), .B0(n8391), .Y(n6120) );
  OAI21XL U15315 ( .A0(n5316), .A1(n6725), .B0(n8391), .Y(n6121) );
  OAI21XL U15316 ( .A0(n5356), .A1(n7673), .B0(n8389), .Y(n6161) );
  OAI21XL U15317 ( .A0(n5357), .A1(n7673), .B0(n8389), .Y(n6162) );
  OAI21XL U15318 ( .A0(n5358), .A1(n7673), .B0(n8389), .Y(n6163) );
  OAI21XL U15319 ( .A0(n5359), .A1(n7673), .B0(n8389), .Y(n6164) );
  OAI21XL U15320 ( .A0(n5360), .A1(n7673), .B0(n8389), .Y(n6165) );
  OAI21XL U15321 ( .A0(n5361), .A1(n6726), .B0(n8389), .Y(n6166) );
  OAI21XL U15322 ( .A0(n5362), .A1(n6726), .B0(n8389), .Y(n6167) );
  OAI21XL U15323 ( .A0(n5363), .A1(n6726), .B0(n8389), .Y(n6168) );
  OAI21XL U15324 ( .A0(n5364), .A1(n6726), .B0(n8389), .Y(n6169) );
  OAI21XL U15325 ( .A0(n5404), .A1(n7674), .B0(n8387), .Y(n6209) );
  OAI21XL U15326 ( .A0(n5405), .A1(n7674), .B0(n8387), .Y(n6210) );
  OAI21XL U15327 ( .A0(n5406), .A1(n7674), .B0(n8387), .Y(n6211) );
  OAI21XL U15328 ( .A0(n5407), .A1(n7674), .B0(n8387), .Y(n6212) );
  OAI21XL U15329 ( .A0(n5408), .A1(n7675), .B0(n8387), .Y(n6213) );
  OAI21XL U15330 ( .A0(n5409), .A1(n7675), .B0(n8387), .Y(n6214) );
  OAI21XL U15331 ( .A0(n5410), .A1(n7675), .B0(n8387), .Y(n6215) );
  OAI21XL U15332 ( .A0(n5411), .A1(n7675), .B0(n8387), .Y(n6216) );
  OAI21XL U15333 ( .A0(n5412), .A1(n7675), .B0(n8387), .Y(n6217) );
  OAI21XL U15334 ( .A0(n5452), .A1(n7677), .B0(n8385), .Y(n6257) );
  OAI21XL U15335 ( .A0(n5453), .A1(n7677), .B0(n8385), .Y(n6258) );
  OAI21XL U15336 ( .A0(n5454), .A1(n7677), .B0(n8385), .Y(n6259) );
  OAI21XL U15337 ( .A0(n5455), .A1(n7677), .B0(n8385), .Y(n6260) );
  OAI21XL U15338 ( .A0(n5456), .A1(n7677), .B0(n8385), .Y(n6261) );
  OAI21XL U15339 ( .A0(n5457), .A1(n6728), .B0(n8385), .Y(n6262) );
  OAI21XL U15340 ( .A0(n5458), .A1(n6728), .B0(n8385), .Y(n6263) );
  OAI21XL U15341 ( .A0(n5459), .A1(n6728), .B0(n8385), .Y(n6264) );
  OAI21XL U15342 ( .A0(n5460), .A1(n6728), .B0(n8385), .Y(n6265) );
  OAI21XL U15343 ( .A0(n5500), .A1(n7678), .B0(n8383), .Y(n6305) );
  OAI21XL U15344 ( .A0(n5501), .A1(n7678), .B0(n8383), .Y(n6306) );
  OAI21XL U15345 ( .A0(n5502), .A1(n7678), .B0(n8383), .Y(n6307) );
  OAI21XL U15346 ( .A0(n5503), .A1(n7679), .B0(n8383), .Y(n6308) );
  OAI21XL U15347 ( .A0(n5504), .A1(n7679), .B0(n8383), .Y(n6309) );
  OAI21XL U15348 ( .A0(n5505), .A1(n7679), .B0(n8383), .Y(n6310) );
  OAI21XL U15349 ( .A0(n5506), .A1(n7679), .B0(n8383), .Y(n6311) );
  OAI21XL U15350 ( .A0(n5507), .A1(n7679), .B0(n8383), .Y(n6312) );
  OAI21XL U15351 ( .A0(n5508), .A1(n7679), .B0(n8383), .Y(n6313) );
  OAI21XL U15352 ( .A0(n5548), .A1(n7681), .B0(n8381), .Y(n6353) );
  OAI21XL U15353 ( .A0(n5549), .A1(n7681), .B0(n8381), .Y(n6354) );
  OAI21XL U15354 ( .A0(n5550), .A1(n7681), .B0(n8381), .Y(n6355) );
  OAI21XL U15355 ( .A0(n5551), .A1(n7681), .B0(n8381), .Y(n6356) );
  OAI21XL U15356 ( .A0(n5552), .A1(n7681), .B0(n8381), .Y(n6357) );
  OAI21XL U15357 ( .A0(n5553), .A1(n6730), .B0(n8381), .Y(n6358) );
  OAI21XL U15358 ( .A0(n5554), .A1(n6730), .B0(n8381), .Y(n6359) );
  OAI21XL U15359 ( .A0(n5555), .A1(n6730), .B0(n8381), .Y(n6360) );
  OAI21XL U15360 ( .A0(n5556), .A1(n6730), .B0(n8381), .Y(n6361) );
  OAI21XL U15361 ( .A0(n5596), .A1(n7683), .B0(n8379), .Y(n6401) );
  OAI21XL U15362 ( .A0(n5597), .A1(n7683), .B0(n8379), .Y(n6402) );
  OAI21XL U15363 ( .A0(n5598), .A1(n7683), .B0(n8379), .Y(n6403) );
  OAI21XL U15364 ( .A0(n5599), .A1(n7683), .B0(n8379), .Y(n6404) );
  OAI21XL U15365 ( .A0(n5600), .A1(n7683), .B0(n8379), .Y(n6405) );
  OAI21XL U15366 ( .A0(n5601), .A1(n6731), .B0(n8379), .Y(n6406) );
  OAI21XL U15367 ( .A0(n5602), .A1(n6731), .B0(n8379), .Y(n6407) );
  OAI21XL U15368 ( .A0(n5603), .A1(n6731), .B0(n8379), .Y(n6408) );
  OAI21XL U15369 ( .A0(n5604), .A1(n6731), .B0(n8379), .Y(n6409) );
  OAI21XL U15370 ( .A0(n5644), .A1(n7685), .B0(n8377), .Y(n6449) );
  OAI21XL U15371 ( .A0(n5645), .A1(n7685), .B0(n8377), .Y(n6450) );
  OAI21XL U15372 ( .A0(n5646), .A1(n7685), .B0(n8377), .Y(n6451) );
  OAI21XL U15373 ( .A0(n5647), .A1(n7685), .B0(n8377), .Y(n6452) );
  OAI21XL U15374 ( .A0(n5648), .A1(n7685), .B0(n8377), .Y(n6453) );
  OAI21XL U15375 ( .A0(n5649), .A1(n6732), .B0(n8377), .Y(n6454) );
  OAI21XL U15376 ( .A0(n5650), .A1(n6732), .B0(n8377), .Y(n6455) );
  OAI21XL U15377 ( .A0(n5651), .A1(n6732), .B0(n8377), .Y(n6456) );
  OAI21XL U15378 ( .A0(n5652), .A1(n6732), .B0(n8377), .Y(n6457) );
  OAI21XL U15379 ( .A0(n5692), .A1(n7697), .B0(n8363), .Y(n6497) );
  OAI21XL U15380 ( .A0(n5693), .A1(n7697), .B0(n8363), .Y(n6498) );
  OAI21XL U15381 ( .A0(n5694), .A1(n7697), .B0(n8363), .Y(n6499) );
  OAI21XL U15382 ( .A0(n5695), .A1(n7697), .B0(n8363), .Y(n6500) );
  OAI21XL U15383 ( .A0(n5696), .A1(n7697), .B0(n8363), .Y(n6501) );
  OAI21XL U15384 ( .A0(n5697), .A1(n6733), .B0(n8363), .Y(n6502) );
  OAI21XL U15385 ( .A0(n5698), .A1(n6733), .B0(n8363), .Y(n6503) );
  OAI21XL U15386 ( .A0(n5699), .A1(n6733), .B0(n8363), .Y(n6504) );
  OAI21XL U15387 ( .A0(n5700), .A1(n6733), .B0(n8363), .Y(n6505) );
  OAI21XL U15388 ( .A0(n4949), .A1(n7698), .B0(n8376), .Y(n5754) );
  OAI21XL U15389 ( .A0(n4950), .A1(n7698), .B0(n8375), .Y(n5755) );
  OAI21XL U15390 ( .A0(n4951), .A1(n7698), .B0(n8376), .Y(n5756) );
  OAI21XL U15391 ( .A0(n4952), .A1(n7698), .B0(n8375), .Y(n5757) );
  OAI21XL U15392 ( .A0(n4953), .A1(n7698), .B0(n215), .Y(n5758) );
  OAI21XL U15393 ( .A0(n4954), .A1(n7698), .B0(n215), .Y(n5759) );
  OAI21XL U15394 ( .A0(n4955), .A1(n7698), .B0(n215), .Y(n5760) );
  OAI21XL U15395 ( .A0(n4956), .A1(n7698), .B0(n8376), .Y(n5761) );
  OAI21XL U15396 ( .A0(n4957), .A1(n7698), .B0(n8376), .Y(n5762) );
  OAI21XL U15397 ( .A0(n4958), .A1(n7698), .B0(n8376), .Y(n5763) );
  OAI21XL U15398 ( .A0(n4959), .A1(n7698), .B0(n8376), .Y(n5764) );
  OAI21XL U15399 ( .A0(n4960), .A1(n7698), .B0(n8376), .Y(n5765) );
  OAI21XL U15400 ( .A0(n4961), .A1(n7698), .B0(n8376), .Y(n5766) );
  OAI21XL U15401 ( .A0(n4962), .A1(n7699), .B0(n8376), .Y(n5767) );
  OAI21XL U15402 ( .A0(n4963), .A1(n7699), .B0(n8376), .Y(n5768) );
  OAI21XL U15403 ( .A0(n4964), .A1(n6719), .B0(n8376), .Y(n5769) );
  OAI21XL U15404 ( .A0(n4965), .A1(n6719), .B0(n8376), .Y(n5770) );
  OAI21XL U15405 ( .A0(n4966), .A1(n6719), .B0(n8376), .Y(n5771) );
  OAI21XL U15406 ( .A0(n4967), .A1(n6719), .B0(n8376), .Y(n5772) );
  OAI21XL U15407 ( .A0(n4968), .A1(n7699), .B0(n8376), .Y(n5773) );
  OAI21XL U15408 ( .A0(n4969), .A1(n7698), .B0(n8375), .Y(n5774) );
  OAI21XL U15409 ( .A0(n4970), .A1(n7698), .B0(n8375), .Y(n5775) );
  OAI21XL U15410 ( .A0(n4971), .A1(n7698), .B0(n8375), .Y(n5776) );
  OAI21XL U15411 ( .A0(n4981), .A1(n7698), .B0(n8375), .Y(n5786) );
  OAI21XL U15412 ( .A0(n4997), .A1(n6720), .B0(n8374), .Y(n5802) );
  OAI21XL U15413 ( .A0(n4998), .A1(n6720), .B0(n8373), .Y(n5803) );
  OAI21XL U15414 ( .A0(n4999), .A1(n6720), .B0(n218), .Y(n5804) );
  OAI21XL U15415 ( .A0(n5000), .A1(n6720), .B0(n218), .Y(n5805) );
  OAI21XL U15416 ( .A0(n5001), .A1(n6720), .B0(n218), .Y(n5806) );
  OAI21XL U15417 ( .A0(n5002), .A1(n7686), .B0(n218), .Y(n5807) );
  OAI21XL U15418 ( .A0(n5003), .A1(n7686), .B0(n218), .Y(n5808) );
  OAI21XL U15419 ( .A0(n5004), .A1(n7686), .B0(n8374), .Y(n5809) );
  OAI21XL U15420 ( .A0(n5005), .A1(n6720), .B0(n8374), .Y(n5810) );
  OAI21XL U15421 ( .A0(n5006), .A1(n6720), .B0(n8374), .Y(n5811) );
  OAI21XL U15422 ( .A0(n5007), .A1(n7686), .B0(n8374), .Y(n5812) );
  OAI21XL U15423 ( .A0(n5008), .A1(n7686), .B0(n8374), .Y(n5813) );
  OAI21XL U15424 ( .A0(n5009), .A1(n7686), .B0(n8374), .Y(n5814) );
  OAI21XL U15425 ( .A0(n5010), .A1(n7686), .B0(n8374), .Y(n5815) );
  OAI21XL U15426 ( .A0(n5011), .A1(n7686), .B0(n8374), .Y(n5816) );
  OAI21XL U15427 ( .A0(n5012), .A1(n7686), .B0(n8374), .Y(n5817) );
  OAI21XL U15428 ( .A0(n5013), .A1(n7686), .B0(n8374), .Y(n5818) );
  OAI21XL U15429 ( .A0(n5014), .A1(n7686), .B0(n8374), .Y(n5819) );
  OAI21XL U15430 ( .A0(n5015), .A1(n7686), .B0(n8374), .Y(n5820) );
  OAI21XL U15431 ( .A0(n5016), .A1(n7686), .B0(n8374), .Y(n5821) );
  OAI21XL U15432 ( .A0(n5017), .A1(n7687), .B0(n8373), .Y(n5822) );
  OAI21XL U15433 ( .A0(n5018), .A1(n7686), .B0(n8373), .Y(n5823) );
  OAI21XL U15434 ( .A0(n5019), .A1(n7686), .B0(n8373), .Y(n5824) );
  OAI21XL U15435 ( .A0(n5029), .A1(n7686), .B0(n8373), .Y(n5834) );
  OAI21XL U15436 ( .A0(n5045), .A1(n7688), .B0(n8372), .Y(n5850) );
  OAI21XL U15437 ( .A0(n5046), .A1(n7688), .B0(n8371), .Y(n5851) );
  OAI21XL U15438 ( .A0(n5047), .A1(n7688), .B0(n222), .Y(n5852) );
  OAI21XL U15439 ( .A0(n5048), .A1(n7688), .B0(n222), .Y(n5853) );
  OAI21XL U15440 ( .A0(n5049), .A1(n7688), .B0(n222), .Y(n5854) );
  OAI21XL U15441 ( .A0(n5050), .A1(n7688), .B0(n222), .Y(n5855) );
  OAI21XL U15442 ( .A0(n5051), .A1(n7688), .B0(n222), .Y(n5856) );
  OAI21XL U15443 ( .A0(n5052), .A1(n7688), .B0(n8372), .Y(n5857) );
  OAI21XL U15444 ( .A0(n5053), .A1(n7688), .B0(n8372), .Y(n5858) );
  OAI21XL U15445 ( .A0(n5054), .A1(n7688), .B0(n8372), .Y(n5859) );
  OAI21XL U15446 ( .A0(n5055), .A1(n7688), .B0(n8372), .Y(n5860) );
  OAI21XL U15447 ( .A0(n5056), .A1(n7688), .B0(n8372), .Y(n5861) );
  OAI21XL U15448 ( .A0(n5057), .A1(n7688), .B0(n8372), .Y(n5862) );
  OAI21XL U15449 ( .A0(n5058), .A1(n7689), .B0(n8372), .Y(n5863) );
  OAI21XL U15450 ( .A0(n5059), .A1(n7689), .B0(n8372), .Y(n5864) );
  OAI21XL U15451 ( .A0(n5060), .A1(n6721), .B0(n8372), .Y(n5865) );
  OAI21XL U15452 ( .A0(n5061), .A1(n6721), .B0(n8372), .Y(n5866) );
  OAI21XL U15453 ( .A0(n5062), .A1(n6721), .B0(n8372), .Y(n5867) );
  OAI21XL U15454 ( .A0(n5063), .A1(n6721), .B0(n8372), .Y(n5868) );
  OAI21XL U15455 ( .A0(n5064), .A1(n7689), .B0(n8372), .Y(n5869) );
  OAI21XL U15456 ( .A0(n5065), .A1(n7688), .B0(n8371), .Y(n5870) );
  OAI21XL U15457 ( .A0(n5066), .A1(n7688), .B0(n8371), .Y(n5871) );
  OAI21XL U15458 ( .A0(n5067), .A1(n7688), .B0(n8371), .Y(n5872) );
  OAI21XL U15459 ( .A0(n5077), .A1(n7688), .B0(n8371), .Y(n5882) );
  OAI21XL U15460 ( .A0(n5093), .A1(n6722), .B0(n8370), .Y(n5898) );
  OAI21XL U15461 ( .A0(n5094), .A1(n6722), .B0(n8369), .Y(n5899) );
  OAI21XL U15462 ( .A0(n5095), .A1(n6722), .B0(n226), .Y(n5900) );
  OAI21XL U15463 ( .A0(n5096), .A1(n6722), .B0(n226), .Y(n5901) );
  OAI21XL U15464 ( .A0(n5097), .A1(n7690), .B0(n226), .Y(n5902) );
  OAI21XL U15465 ( .A0(n5098), .A1(n7690), .B0(n226), .Y(n5903) );
  OAI21XL U15466 ( .A0(n5099), .A1(n7690), .B0(n226), .Y(n5904) );
  OAI21XL U15467 ( .A0(n5100), .A1(n6722), .B0(n8370), .Y(n5905) );
  OAI21XL U15468 ( .A0(n5101), .A1(n6722), .B0(n8370), .Y(n5906) );
  OAI21XL U15469 ( .A0(n5102), .A1(n7690), .B0(n8370), .Y(n5907) );
  OAI21XL U15470 ( .A0(n5103), .A1(n7690), .B0(n8370), .Y(n5908) );
  OAI21XL U15471 ( .A0(n5104), .A1(n7690), .B0(n8370), .Y(n5909) );
  OAI21XL U15472 ( .A0(n5105), .A1(n7690), .B0(n8370), .Y(n5910) );
  OAI21XL U15473 ( .A0(n5106), .A1(n7690), .B0(n8370), .Y(n5911) );
  OAI21XL U15474 ( .A0(n5107), .A1(n7690), .B0(n8370), .Y(n5912) );
  OAI21XL U15475 ( .A0(n5108), .A1(n7690), .B0(n8370), .Y(n5913) );
  OAI21XL U15476 ( .A0(n5109), .A1(n7690), .B0(n8370), .Y(n5914) );
  OAI21XL U15477 ( .A0(n5110), .A1(n7690), .B0(n8370), .Y(n5915) );
  OAI21XL U15478 ( .A0(n5111), .A1(n7690), .B0(n8370), .Y(n5916) );
  OAI21XL U15479 ( .A0(n5112), .A1(n7690), .B0(n8370), .Y(n5917) );
  OAI21XL U15480 ( .A0(n5113), .A1(n7690), .B0(n8369), .Y(n5918) );
  OAI21XL U15481 ( .A0(n5114), .A1(n7690), .B0(n8369), .Y(n5919) );
  OAI21XL U15482 ( .A0(n5115), .A1(n7690), .B0(n8369), .Y(n5920) );
  OAI21XL U15483 ( .A0(n5125), .A1(n6722), .B0(n8369), .Y(n5930) );
  OAI21XL U15484 ( .A0(n5141), .A1(n7692), .B0(n8368), .Y(n5946) );
  OAI21XL U15485 ( .A0(n5142), .A1(n7692), .B0(n8367), .Y(n5947) );
  OAI21XL U15486 ( .A0(n5143), .A1(n7692), .B0(n230), .Y(n5948) );
  OAI21XL U15487 ( .A0(n5144), .A1(n7692), .B0(n230), .Y(n5949) );
  OAI21XL U15488 ( .A0(n5145), .A1(n7692), .B0(n230), .Y(n5950) );
  OAI21XL U15489 ( .A0(n5146), .A1(n7692), .B0(n230), .Y(n5951) );
  OAI21XL U15490 ( .A0(n5147), .A1(n7692), .B0(n230), .Y(n5952) );
  OAI21XL U15491 ( .A0(n5148), .A1(n7692), .B0(n8368), .Y(n5953) );
  OAI21XL U15492 ( .A0(n5149), .A1(n7692), .B0(n8368), .Y(n5954) );
  OAI21XL U15493 ( .A0(n5150), .A1(n7692), .B0(n8368), .Y(n5955) );
  OAI21XL U15494 ( .A0(n5151), .A1(n7692), .B0(n8368), .Y(n5956) );
  OAI21XL U15495 ( .A0(n5152), .A1(n7692), .B0(n8368), .Y(n5957) );
  OAI21XL U15496 ( .A0(n5153), .A1(n7692), .B0(n8368), .Y(n5958) );
  OAI21XL U15497 ( .A0(n5154), .A1(n7693), .B0(n8368), .Y(n5959) );
  OAI21XL U15498 ( .A0(n5155), .A1(n7693), .B0(n8368), .Y(n5960) );
  OAI21XL U15499 ( .A0(n5156), .A1(n6723), .B0(n8368), .Y(n5961) );
  OAI21XL U15500 ( .A0(n5157), .A1(n6723), .B0(n8368), .Y(n5962) );
  OAI21XL U15501 ( .A0(n5158), .A1(n6723), .B0(n8368), .Y(n5963) );
  OAI21XL U15502 ( .A0(n5159), .A1(n6723), .B0(n8368), .Y(n5964) );
  OAI21XL U15503 ( .A0(n5160), .A1(n7693), .B0(n8368), .Y(n5965) );
  OAI21XL U15504 ( .A0(n5161), .A1(n7692), .B0(n8367), .Y(n5966) );
  OAI21XL U15505 ( .A0(n5162), .A1(n7692), .B0(n8367), .Y(n5967) );
  OAI21XL U15506 ( .A0(n5163), .A1(n7692), .B0(n8367), .Y(n5968) );
  OAI21XL U15507 ( .A0(n5173), .A1(n7692), .B0(n8367), .Y(n5978) );
  OAI21XL U15508 ( .A0(n5189), .A1(n7694), .B0(n8366), .Y(n5994) );
  OAI21XL U15509 ( .A0(n5190), .A1(n7694), .B0(n8365), .Y(n5995) );
  OAI21XL U15510 ( .A0(n5191), .A1(n7694), .B0(n234), .Y(n5996) );
  OAI21XL U15511 ( .A0(n5192), .A1(n7694), .B0(n234), .Y(n5997) );
  OAI21XL U15512 ( .A0(n5193), .A1(n7694), .B0(n234), .Y(n5998) );
  OAI21XL U15513 ( .A0(n5194), .A1(n7694), .B0(n234), .Y(n5999) );
  OAI21XL U15514 ( .A0(n5195), .A1(n7694), .B0(n234), .Y(n6000) );
  OAI21XL U15515 ( .A0(n5196), .A1(n7694), .B0(n8366), .Y(n6001) );
  OAI21XL U15516 ( .A0(n5197), .A1(n7694), .B0(n8366), .Y(n6002) );
  OAI21XL U15517 ( .A0(n5198), .A1(n7694), .B0(n8366), .Y(n6003) );
  OAI21XL U15518 ( .A0(n5199), .A1(n7694), .B0(n8366), .Y(n6004) );
  OAI21XL U15519 ( .A0(n5200), .A1(n7694), .B0(n8366), .Y(n6005) );
  OAI21XL U15520 ( .A0(n5201), .A1(n7694), .B0(n8366), .Y(n6006) );
  OAI21XL U15521 ( .A0(n5202), .A1(n7695), .B0(n8366), .Y(n6007) );
  OAI21XL U15522 ( .A0(n5203), .A1(n7695), .B0(n8366), .Y(n6008) );
  OAI21XL U15523 ( .A0(n5204), .A1(n6724), .B0(n8366), .Y(n6009) );
  OAI21XL U15524 ( .A0(n5205), .A1(n6724), .B0(n8366), .Y(n6010) );
  OAI21XL U15525 ( .A0(n5206), .A1(n6724), .B0(n8366), .Y(n6011) );
  OAI21XL U15526 ( .A0(n5207), .A1(n6724), .B0(n8366), .Y(n6012) );
  OAI21XL U15527 ( .A0(n5208), .A1(n7695), .B0(n8366), .Y(n6013) );
  OAI21XL U15528 ( .A0(n5209), .A1(n7694), .B0(n8365), .Y(n6014) );
  OAI21XL U15529 ( .A0(n5210), .A1(n7694), .B0(n8365), .Y(n6015) );
  OAI21XL U15530 ( .A0(n5211), .A1(n7694), .B0(n8365), .Y(n6016) );
  OAI21XL U15531 ( .A0(n5221), .A1(n7694), .B0(n8365), .Y(n6026) );
  OAI21XL U15532 ( .A0(n5237), .A1(n7668), .B0(n8394), .Y(n6042) );
  OAI21XL U15533 ( .A0(n5238), .A1(n7668), .B0(n8393), .Y(n6043) );
  OAI21XL U15534 ( .A0(n5239), .A1(n7668), .B0(n164), .Y(n6044) );
  OAI21XL U15535 ( .A0(n5240), .A1(n7668), .B0(n164), .Y(n6045) );
  OAI21XL U15536 ( .A0(n5241), .A1(n7668), .B0(n164), .Y(n6046) );
  OAI21XL U15537 ( .A0(n5242), .A1(n7668), .B0(n164), .Y(n6047) );
  OAI21XL U15538 ( .A0(n5243), .A1(n7668), .B0(n164), .Y(n6048) );
  OAI21XL U15539 ( .A0(n5244), .A1(n7668), .B0(n8394), .Y(n6049) );
  OAI21XL U15540 ( .A0(n5245), .A1(n7668), .B0(n8394), .Y(n6050) );
  OAI21XL U15541 ( .A0(n5246), .A1(n7668), .B0(n8394), .Y(n6051) );
  OAI21XL U15542 ( .A0(n5247), .A1(n7668), .B0(n8394), .Y(n6052) );
  OAI21XL U15543 ( .A0(n5248), .A1(n7668), .B0(n8394), .Y(n6053) );
  OAI21XL U15544 ( .A0(n5249), .A1(n7668), .B0(n8394), .Y(n6054) );
  OAI21XL U15545 ( .A0(n5250), .A1(n7669), .B0(n8394), .Y(n6055) );
  OAI21XL U15546 ( .A0(n5251), .A1(n7669), .B0(n8394), .Y(n6056) );
  OAI21XL U15547 ( .A0(n5252), .A1(n6734), .B0(n8394), .Y(n6057) );
  OAI21XL U15548 ( .A0(n5253), .A1(n6734), .B0(n8394), .Y(n6058) );
  OAI21XL U15549 ( .A0(n5254), .A1(n6734), .B0(n8394), .Y(n6059) );
  OAI21XL U15550 ( .A0(n5255), .A1(n6734), .B0(n8394), .Y(n6060) );
  OAI21XL U15551 ( .A0(n5256), .A1(n7669), .B0(n8394), .Y(n6061) );
  OAI21XL U15552 ( .A0(n5257), .A1(n7668), .B0(n8393), .Y(n6062) );
  OAI21XL U15553 ( .A0(n5258), .A1(n7668), .B0(n8393), .Y(n6063) );
  OAI21XL U15554 ( .A0(n5259), .A1(n7668), .B0(n8393), .Y(n6064) );
  OAI21XL U15555 ( .A0(n5269), .A1(n7668), .B0(n8393), .Y(n6074) );
  OAI21XL U15556 ( .A0(n5285), .A1(n7670), .B0(n8392), .Y(n6090) );
  OAI21XL U15557 ( .A0(n5286), .A1(n7670), .B0(n8391), .Y(n6091) );
  OAI21XL U15558 ( .A0(n5287), .A1(n7670), .B0(n183), .Y(n6092) );
  OAI21XL U15559 ( .A0(n5288), .A1(n7670), .B0(n183), .Y(n6093) );
  OAI21XL U15560 ( .A0(n5289), .A1(n7670), .B0(n183), .Y(n6094) );
  OAI21XL U15561 ( .A0(n5290), .A1(n7670), .B0(n183), .Y(n6095) );
  OAI21XL U15562 ( .A0(n5291), .A1(n7670), .B0(n183), .Y(n6096) );
  OAI21XL U15563 ( .A0(n5292), .A1(n7670), .B0(n8392), .Y(n6097) );
  OAI21XL U15564 ( .A0(n5293), .A1(n7670), .B0(n8392), .Y(n6098) );
  OAI21XL U15565 ( .A0(n5294), .A1(n7670), .B0(n8392), .Y(n6099) );
  OAI21XL U15566 ( .A0(n5295), .A1(n7670), .B0(n8392), .Y(n6100) );
  OAI21XL U15567 ( .A0(n5296), .A1(n7670), .B0(n8392), .Y(n6101) );
  OAI21XL U15568 ( .A0(n5297), .A1(n7670), .B0(n8392), .Y(n6102) );
  OAI21XL U15569 ( .A0(n5298), .A1(n7671), .B0(n8392), .Y(n6103) );
  OAI21XL U15570 ( .A0(n5299), .A1(n7671), .B0(n8392), .Y(n6104) );
  OAI21XL U15571 ( .A0(n5300), .A1(n6725), .B0(n8392), .Y(n6105) );
  OAI21XL U15572 ( .A0(n5301), .A1(n6725), .B0(n8392), .Y(n6106) );
  OAI21XL U15573 ( .A0(n5302), .A1(n6725), .B0(n8392), .Y(n6107) );
  OAI21XL U15574 ( .A0(n5303), .A1(n6725), .B0(n8392), .Y(n6108) );
  OAI21XL U15575 ( .A0(n5304), .A1(n7671), .B0(n8392), .Y(n6109) );
  OAI21XL U15576 ( .A0(n5305), .A1(n7670), .B0(n8391), .Y(n6110) );
  OAI21XL U15577 ( .A0(n5306), .A1(n7670), .B0(n8391), .Y(n6111) );
  OAI21XL U15578 ( .A0(n5307), .A1(n7670), .B0(n8391), .Y(n6112) );
  OAI21XL U15579 ( .A0(n5317), .A1(n7670), .B0(n8391), .Y(n6122) );
  OAI21XL U15580 ( .A0(n5333), .A1(n7672), .B0(n8390), .Y(n6138) );
  OAI21XL U15581 ( .A0(n5334), .A1(n7672), .B0(n8389), .Y(n6139) );
  OAI21XL U15582 ( .A0(n5335), .A1(n7672), .B0(n187), .Y(n6140) );
  OAI21XL U15583 ( .A0(n5336), .A1(n7672), .B0(n187), .Y(n6141) );
  OAI21XL U15584 ( .A0(n5337), .A1(n7672), .B0(n187), .Y(n6142) );
  OAI21XL U15585 ( .A0(n5338), .A1(n7672), .B0(n187), .Y(n6143) );
  OAI21XL U15586 ( .A0(n5339), .A1(n7672), .B0(n187), .Y(n6144) );
  OAI21XL U15587 ( .A0(n5340), .A1(n7672), .B0(n8390), .Y(n6145) );
  OAI21XL U15588 ( .A0(n5341), .A1(n7672), .B0(n8390), .Y(n6146) );
  OAI21XL U15589 ( .A0(n5342), .A1(n7672), .B0(n8390), .Y(n6147) );
  OAI21XL U15590 ( .A0(n5343), .A1(n7672), .B0(n8390), .Y(n6148) );
  OAI21XL U15591 ( .A0(n5344), .A1(n7672), .B0(n8390), .Y(n6149) );
  OAI21XL U15592 ( .A0(n5345), .A1(n7672), .B0(n8390), .Y(n6150) );
  OAI21XL U15593 ( .A0(n5346), .A1(n7673), .B0(n8390), .Y(n6151) );
  OAI21XL U15594 ( .A0(n5347), .A1(n7673), .B0(n8390), .Y(n6152) );
  OAI21XL U15595 ( .A0(n5348), .A1(n6726), .B0(n8390), .Y(n6153) );
  OAI21XL U15596 ( .A0(n5349), .A1(n6726), .B0(n8390), .Y(n6154) );
  OAI21XL U15597 ( .A0(n5350), .A1(n6726), .B0(n8390), .Y(n6155) );
  OAI21XL U15598 ( .A0(n5351), .A1(n6726), .B0(n8390), .Y(n6156) );
  OAI21XL U15599 ( .A0(n5352), .A1(n7673), .B0(n8390), .Y(n6157) );
  OAI21XL U15600 ( .A0(n5353), .A1(n7672), .B0(n8389), .Y(n6158) );
  OAI21XL U15601 ( .A0(n5354), .A1(n7672), .B0(n8389), .Y(n6159) );
  OAI21XL U15602 ( .A0(n5355), .A1(n7672), .B0(n8389), .Y(n6160) );
  OAI21XL U15603 ( .A0(n5365), .A1(n7672), .B0(n8389), .Y(n6170) );
  OAI21XL U15604 ( .A0(n5381), .A1(n6727), .B0(n8388), .Y(n6186) );
  OAI21XL U15605 ( .A0(n5382), .A1(n6727), .B0(n8387), .Y(n6187) );
  OAI21XL U15606 ( .A0(n5383), .A1(n6727), .B0(n191), .Y(n6188) );
  OAI21XL U15607 ( .A0(n5384), .A1(n6727), .B0(n191), .Y(n6189) );
  OAI21XL U15608 ( .A0(n5385), .A1(n6727), .B0(n191), .Y(n6190) );
  OAI21XL U15609 ( .A0(n5386), .A1(n7674), .B0(n191), .Y(n6191) );
  OAI21XL U15610 ( .A0(n5387), .A1(n7674), .B0(n191), .Y(n6192) );
  OAI21XL U15611 ( .A0(n5388), .A1(n7674), .B0(n8388), .Y(n6193) );
  OAI21XL U15612 ( .A0(n5389), .A1(n6727), .B0(n8388), .Y(n6194) );
  OAI21XL U15613 ( .A0(n5390), .A1(n6727), .B0(n8388), .Y(n6195) );
  OAI21XL U15614 ( .A0(n5391), .A1(n7674), .B0(n8388), .Y(n6196) );
  OAI21XL U15615 ( .A0(n5392), .A1(n7674), .B0(n8388), .Y(n6197) );
  OAI21XL U15616 ( .A0(n5393), .A1(n7674), .B0(n8388), .Y(n6198) );
  OAI21XL U15617 ( .A0(n5394), .A1(n7674), .B0(n8388), .Y(n6199) );
  OAI21XL U15618 ( .A0(n5395), .A1(n7674), .B0(n8388), .Y(n6200) );
  OAI21XL U15619 ( .A0(n5396), .A1(n7674), .B0(n8388), .Y(n6201) );
  OAI21XL U15620 ( .A0(n5397), .A1(n7674), .B0(n8388), .Y(n6202) );
  OAI21XL U15621 ( .A0(n5398), .A1(n7674), .B0(n8388), .Y(n6203) );
  OAI21XL U15622 ( .A0(n5399), .A1(n7674), .B0(n8388), .Y(n6204) );
  OAI21XL U15623 ( .A0(n5400), .A1(n7674), .B0(n8388), .Y(n6205) );
  OAI21XL U15624 ( .A0(n5401), .A1(n7675), .B0(n8387), .Y(n6206) );
  OAI21XL U15625 ( .A0(n5402), .A1(n7674), .B0(n8387), .Y(n6207) );
  OAI21XL U15626 ( .A0(n5403), .A1(n7674), .B0(n8387), .Y(n6208) );
  OAI21XL U15627 ( .A0(n5413), .A1(n7674), .B0(n8387), .Y(n6218) );
  OAI21XL U15628 ( .A0(n5429), .A1(n7676), .B0(n8386), .Y(n6234) );
  OAI21XL U15629 ( .A0(n5430), .A1(n7676), .B0(n8385), .Y(n6235) );
  OAI21XL U15630 ( .A0(n5431), .A1(n7676), .B0(n8386), .Y(n6236) );
  OAI21XL U15631 ( .A0(n5432), .A1(n7676), .B0(n8385), .Y(n6237) );
  OAI21XL U15632 ( .A0(n5433), .A1(n7676), .B0(n195), .Y(n6238) );
  OAI21XL U15633 ( .A0(n5434), .A1(n7676), .B0(n195), .Y(n6239) );
  OAI21XL U15634 ( .A0(n5435), .A1(n7676), .B0(n195), .Y(n6240) );
  OAI21XL U15635 ( .A0(n5436), .A1(n7676), .B0(n8386), .Y(n6241) );
  OAI21XL U15636 ( .A0(n5437), .A1(n7676), .B0(n8386), .Y(n6242) );
  OAI21XL U15637 ( .A0(n5438), .A1(n7676), .B0(n8386), .Y(n6243) );
  OAI21XL U15638 ( .A0(n5439), .A1(n7676), .B0(n8386), .Y(n6244) );
  OAI21XL U15639 ( .A0(n5440), .A1(n7676), .B0(n8386), .Y(n6245) );
  OAI21XL U15640 ( .A0(n5441), .A1(n7676), .B0(n8386), .Y(n6246) );
  OAI21XL U15641 ( .A0(n5442), .A1(n7677), .B0(n8386), .Y(n6247) );
  OAI21XL U15642 ( .A0(n5443), .A1(n7677), .B0(n8386), .Y(n6248) );
  OAI21XL U15643 ( .A0(n5444), .A1(n6728), .B0(n8386), .Y(n6249) );
  OAI21XL U15644 ( .A0(n5445), .A1(n6728), .B0(n8386), .Y(n6250) );
  OAI21XL U15645 ( .A0(n5446), .A1(n6728), .B0(n8386), .Y(n6251) );
  OAI21XL U15646 ( .A0(n5447), .A1(n6728), .B0(n8386), .Y(n6252) );
  OAI21XL U15647 ( .A0(n5448), .A1(n7677), .B0(n8386), .Y(n6253) );
  OAI21XL U15648 ( .A0(n5449), .A1(n7676), .B0(n8385), .Y(n6254) );
  OAI21XL U15649 ( .A0(n5450), .A1(n7676), .B0(n8385), .Y(n6255) );
  OAI21XL U15650 ( .A0(n5451), .A1(n7676), .B0(n8385), .Y(n6256) );
  OAI21XL U15651 ( .A0(n5461), .A1(n7676), .B0(n8385), .Y(n6266) );
  OAI21XL U15652 ( .A0(n5477), .A1(n6729), .B0(n8384), .Y(n6282) );
  OAI21XL U15653 ( .A0(n5478), .A1(n6729), .B0(n8383), .Y(n6283) );
  OAI21XL U15654 ( .A0(n5479), .A1(n6729), .B0(n199), .Y(n6284) );
  OAI21XL U15655 ( .A0(n5480), .A1(n6729), .B0(n199), .Y(n6285) );
  OAI21XL U15656 ( .A0(n5481), .A1(n7678), .B0(n199), .Y(n6286) );
  OAI21XL U15657 ( .A0(n5482), .A1(n7678), .B0(n199), .Y(n6287) );
  OAI21XL U15658 ( .A0(n5483), .A1(n7678), .B0(n199), .Y(n6288) );
  OAI21XL U15659 ( .A0(n5484), .A1(n6729), .B0(n8384), .Y(n6289) );
  OAI21XL U15660 ( .A0(n5485), .A1(n6729), .B0(n8384), .Y(n6290) );
  OAI21XL U15661 ( .A0(n5486), .A1(n7678), .B0(n8384), .Y(n6291) );
  OAI21XL U15662 ( .A0(n5487), .A1(n7678), .B0(n8384), .Y(n6292) );
  OAI21XL U15663 ( .A0(n5488), .A1(n7678), .B0(n8384), .Y(n6293) );
  OAI21XL U15664 ( .A0(n5489), .A1(n7678), .B0(n8384), .Y(n6294) );
  OAI21XL U15665 ( .A0(n5490), .A1(n7678), .B0(n8384), .Y(n6295) );
  OAI21XL U15666 ( .A0(n5491), .A1(n7678), .B0(n8384), .Y(n6296) );
  OAI21XL U15667 ( .A0(n5492), .A1(n7678), .B0(n8384), .Y(n6297) );
  OAI21XL U15668 ( .A0(n5493), .A1(n7678), .B0(n8384), .Y(n6298) );
  OAI21XL U15669 ( .A0(n5494), .A1(n7678), .B0(n8384), .Y(n6299) );
  OAI21XL U15670 ( .A0(n5495), .A1(n7678), .B0(n8384), .Y(n6300) );
  OAI21XL U15671 ( .A0(n5496), .A1(n7678), .B0(n8384), .Y(n6301) );
  OAI21XL U15672 ( .A0(n5497), .A1(n7678), .B0(n8383), .Y(n6302) );
  OAI21XL U15673 ( .A0(n5498), .A1(n7678), .B0(n8383), .Y(n6303) );
  OAI21XL U15674 ( .A0(n5499), .A1(n7678), .B0(n8383), .Y(n6304) );
  OAI21XL U15675 ( .A0(n5509), .A1(n6729), .B0(n8383), .Y(n6314) );
  OAI21XL U15676 ( .A0(n5525), .A1(n7680), .B0(n8382), .Y(n6330) );
  OAI21XL U15677 ( .A0(n5526), .A1(n7680), .B0(n8381), .Y(n6331) );
  OAI21XL U15678 ( .A0(n5527), .A1(n7680), .B0(n203), .Y(n6332) );
  OAI21XL U15679 ( .A0(n5528), .A1(n7680), .B0(n203), .Y(n6333) );
  OAI21XL U15680 ( .A0(n5529), .A1(n7680), .B0(n203), .Y(n6334) );
  OAI21XL U15681 ( .A0(n5530), .A1(n7680), .B0(n203), .Y(n6335) );
  OAI21XL U15682 ( .A0(n5531), .A1(n7680), .B0(n203), .Y(n6336) );
  OAI21XL U15683 ( .A0(n5532), .A1(n7680), .B0(n8382), .Y(n6337) );
  OAI21XL U15684 ( .A0(n5533), .A1(n7680), .B0(n8382), .Y(n6338) );
  OAI21XL U15685 ( .A0(n5534), .A1(n7680), .B0(n8382), .Y(n6339) );
  OAI21XL U15686 ( .A0(n5535), .A1(n7680), .B0(n8382), .Y(n6340) );
  OAI21XL U15687 ( .A0(n5536), .A1(n7680), .B0(n8382), .Y(n6341) );
  OAI21XL U15688 ( .A0(n5537), .A1(n7680), .B0(n8382), .Y(n6342) );
  OAI21XL U15689 ( .A0(n5538), .A1(n7681), .B0(n8382), .Y(n6343) );
  OAI21XL U15690 ( .A0(n5539), .A1(n7681), .B0(n8382), .Y(n6344) );
  OAI21XL U15691 ( .A0(n5540), .A1(n6730), .B0(n8382), .Y(n6345) );
  OAI21XL U15692 ( .A0(n5541), .A1(n6730), .B0(n8382), .Y(n6346) );
  OAI21XL U15693 ( .A0(n5542), .A1(n6730), .B0(n8382), .Y(n6347) );
  OAI21XL U15694 ( .A0(n5543), .A1(n6730), .B0(n8382), .Y(n6348) );
  OAI21XL U15695 ( .A0(n5544), .A1(n7681), .B0(n8382), .Y(n6349) );
  OAI21XL U15696 ( .A0(n5545), .A1(n7680), .B0(n8381), .Y(n6350) );
  OAI21XL U15697 ( .A0(n5546), .A1(n7680), .B0(n8381), .Y(n6351) );
  OAI21XL U15698 ( .A0(n5547), .A1(n7680), .B0(n8381), .Y(n6352) );
  OAI21XL U15699 ( .A0(n5557), .A1(n7680), .B0(n8381), .Y(n6362) );
  OAI21XL U15700 ( .A0(n5573), .A1(n7682), .B0(n8380), .Y(n6378) );
  OAI21XL U15701 ( .A0(n5574), .A1(n7682), .B0(n8379), .Y(n6379) );
  OAI21XL U15702 ( .A0(n5575), .A1(n7682), .B0(n207), .Y(n6380) );
  OAI21XL U15703 ( .A0(n5576), .A1(n7682), .B0(n207), .Y(n6381) );
  OAI21XL U15704 ( .A0(n5577), .A1(n7682), .B0(n207), .Y(n6382) );
  OAI21XL U15705 ( .A0(n5578), .A1(n7682), .B0(n207), .Y(n6383) );
  OAI21XL U15706 ( .A0(n5579), .A1(n7682), .B0(n207), .Y(n6384) );
  OAI21XL U15707 ( .A0(n5580), .A1(n7682), .B0(n8380), .Y(n6385) );
  OAI21XL U15708 ( .A0(n5581), .A1(n7682), .B0(n8380), .Y(n6386) );
  OAI21XL U15709 ( .A0(n5582), .A1(n7682), .B0(n8380), .Y(n6387) );
  OAI21XL U15710 ( .A0(n5583), .A1(n7682), .B0(n8380), .Y(n6388) );
  OAI21XL U15711 ( .A0(n5584), .A1(n7682), .B0(n8380), .Y(n6389) );
  OAI21XL U15712 ( .A0(n5585), .A1(n7682), .B0(n8380), .Y(n6390) );
  OAI21XL U15713 ( .A0(n5586), .A1(n7683), .B0(n8380), .Y(n6391) );
  OAI21XL U15714 ( .A0(n5587), .A1(n7683), .B0(n8380), .Y(n6392) );
  OAI21XL U15715 ( .A0(n5588), .A1(n6731), .B0(n8380), .Y(n6393) );
  OAI21XL U15716 ( .A0(n5589), .A1(n6731), .B0(n8380), .Y(n6394) );
  OAI21XL U15717 ( .A0(n5590), .A1(n6731), .B0(n8380), .Y(n6395) );
  OAI21XL U15718 ( .A0(n5591), .A1(n6731), .B0(n8380), .Y(n6396) );
  OAI21XL U15719 ( .A0(n5592), .A1(n7683), .B0(n8380), .Y(n6397) );
  OAI21XL U15720 ( .A0(n5593), .A1(n7682), .B0(n8379), .Y(n6398) );
  OAI21XL U15721 ( .A0(n5594), .A1(n7682), .B0(n8379), .Y(n6399) );
  OAI21XL U15722 ( .A0(n5595), .A1(n7682), .B0(n8379), .Y(n6400) );
  OAI21XL U15723 ( .A0(n5605), .A1(n7682), .B0(n8379), .Y(n6410) );
  OAI21XL U15724 ( .A0(n5621), .A1(n7684), .B0(n8378), .Y(n6426) );
  OAI21XL U15725 ( .A0(n5622), .A1(n7684), .B0(n8377), .Y(n6427) );
  OAI21XL U15726 ( .A0(n5623), .A1(n7684), .B0(n8378), .Y(n6428) );
  OAI21XL U15727 ( .A0(n5624), .A1(n7684), .B0(n8377), .Y(n6429) );
  OAI21XL U15728 ( .A0(n5625), .A1(n7684), .B0(n211), .Y(n6430) );
  OAI21XL U15729 ( .A0(n5626), .A1(n7684), .B0(n211), .Y(n6431) );
  OAI21XL U15730 ( .A0(n5627), .A1(n7684), .B0(n211), .Y(n6432) );
  OAI21XL U15731 ( .A0(n5628), .A1(n7684), .B0(n8378), .Y(n6433) );
  OAI21XL U15732 ( .A0(n5629), .A1(n7684), .B0(n8378), .Y(n6434) );
  OAI21XL U15733 ( .A0(n5630), .A1(n7684), .B0(n8378), .Y(n6435) );
  OAI21XL U15734 ( .A0(n5631), .A1(n7684), .B0(n8378), .Y(n6436) );
  OAI21XL U15735 ( .A0(n5632), .A1(n7684), .B0(n8378), .Y(n6437) );
  OAI21XL U15736 ( .A0(n5633), .A1(n7684), .B0(n8378), .Y(n6438) );
  OAI21XL U15737 ( .A0(n5634), .A1(n7685), .B0(n8378), .Y(n6439) );
  OAI21XL U15738 ( .A0(n5635), .A1(n7685), .B0(n8378), .Y(n6440) );
  OAI21XL U15739 ( .A0(n5636), .A1(n6732), .B0(n8378), .Y(n6441) );
  OAI21XL U15740 ( .A0(n5637), .A1(n6732), .B0(n8378), .Y(n6442) );
  OAI21XL U15741 ( .A0(n5638), .A1(n6732), .B0(n8378), .Y(n6443) );
  OAI21XL U15742 ( .A0(n5639), .A1(n6732), .B0(n8378), .Y(n6444) );
  OAI21XL U15743 ( .A0(n5640), .A1(n7685), .B0(n8378), .Y(n6445) );
  OAI21XL U15744 ( .A0(n5641), .A1(n7684), .B0(n8377), .Y(n6446) );
  OAI21XL U15745 ( .A0(n5642), .A1(n7684), .B0(n8377), .Y(n6447) );
  OAI21XL U15746 ( .A0(n5643), .A1(n7684), .B0(n8377), .Y(n6448) );
  OAI21XL U15747 ( .A0(n5653), .A1(n7684), .B0(n8377), .Y(n6458) );
  OAI21XL U15748 ( .A0(n5669), .A1(n7696), .B0(n8364), .Y(n6474) );
  OAI21XL U15749 ( .A0(n5670), .A1(n7696), .B0(n8363), .Y(n6475) );
  OAI21XL U15750 ( .A0(n5671), .A1(n7696), .B0(n238), .Y(n6476) );
  OAI21XL U15751 ( .A0(n5672), .A1(n7696), .B0(n238), .Y(n6477) );
  OAI21XL U15752 ( .A0(n5673), .A1(n7696), .B0(n238), .Y(n6478) );
  OAI21XL U15753 ( .A0(n5674), .A1(n7696), .B0(n238), .Y(n6479) );
  OAI21XL U15754 ( .A0(n5675), .A1(n7696), .B0(n238), .Y(n6480) );
  OAI21XL U15755 ( .A0(n5676), .A1(n7696), .B0(n8364), .Y(n6481) );
  OAI21XL U15756 ( .A0(n5677), .A1(n7696), .B0(n8364), .Y(n6482) );
  OAI21XL U15757 ( .A0(n5678), .A1(n7696), .B0(n8364), .Y(n6483) );
  OAI21XL U15758 ( .A0(n5679), .A1(n7696), .B0(n8364), .Y(n6484) );
  OAI21XL U15759 ( .A0(n5680), .A1(n7696), .B0(n8364), .Y(n6485) );
  OAI21XL U15760 ( .A0(n5681), .A1(n7696), .B0(n8364), .Y(n6486) );
  OAI21XL U15761 ( .A0(n5682), .A1(n7697), .B0(n8364), .Y(n6487) );
  OAI21XL U15762 ( .A0(n5683), .A1(n7697), .B0(n8364), .Y(n6488) );
  OAI21XL U15763 ( .A0(n5684), .A1(n6733), .B0(n8364), .Y(n6489) );
  OAI21XL U15764 ( .A0(n5685), .A1(n6733), .B0(n8364), .Y(n6490) );
  OAI21XL U15765 ( .A0(n5686), .A1(n6733), .B0(n8364), .Y(n6491) );
  OAI21XL U15766 ( .A0(n5687), .A1(n6733), .B0(n8364), .Y(n6492) );
  OAI21XL U15767 ( .A0(n5688), .A1(n7697), .B0(n8364), .Y(n6493) );
  OAI21XL U15768 ( .A0(n5689), .A1(n7696), .B0(n8363), .Y(n6494) );
  OAI21XL U15769 ( .A0(n5690), .A1(n7696), .B0(n8363), .Y(n6495) );
  OAI21XL U15770 ( .A0(n5691), .A1(n7696), .B0(n8363), .Y(n6496) );
  OAI21XL U15771 ( .A0(n5704), .A1(n7696), .B0(n8363), .Y(n6506) );
  NAND4X1 U15772 ( .A(n84), .B(n83), .C(n82), .D(n81), .Y(n4889) );
  NAND4X1 U15773 ( .A(n91), .B(n90), .C(n89), .D(n88), .Y(n4890) );
  NAND4X1 U15774 ( .A(n98), .B(n97), .C(n96), .D(n95), .Y(n4891) );
  AND2X2 U15775 ( .A(n74), .B(n3148), .Y(n3078) );
  NOR2BX1 U15776 ( .AN(N35084), .B(n8398), .Y(outCount_next[0]) );
  AND2X2 U15777 ( .A(N34939), .B(N35192), .Y(N34944) );
  MX4X1 U15778 ( .A(n7239), .B(n7237), .C(n7238), .D(n7236), .S0(n7356), .S1(
        n7359), .Y(N34939) );
  AND2X2 U15779 ( .A(N34938), .B(N35192), .Y(N34945) );
  MX4X1 U15780 ( .A(n7243), .B(n7241), .C(n7242), .D(n7240), .S0(n7356), .S1(
        n7360), .Y(N34938) );
  AND2X2 U15781 ( .A(N34937), .B(N35192), .Y(N34946) );
  MX4X1 U15782 ( .A(n7247), .B(n7245), .C(n7246), .D(n7244), .S0(n7356), .S1(
        n7359), .Y(N34937) );
  AND2X2 U15783 ( .A(N34936), .B(N35192), .Y(N34947) );
  MX4X1 U15784 ( .A(n7251), .B(n7249), .C(n7250), .D(n7248), .S0(n7356), .S1(
        n7360), .Y(N34936) );
  AND2X2 U15785 ( .A(N34935), .B(N35192), .Y(N34948) );
  MX4X1 U15786 ( .A(n7255), .B(n7253), .C(n7254), .D(n7252), .S0(n7357), .S1(
        n7359), .Y(N34935) );
  AND2X2 U15787 ( .A(N34934), .B(N35192), .Y(N34949) );
  MX4X1 U15788 ( .A(n7259), .B(n7257), .C(n7258), .D(n7256), .S0(n7357), .S1(
        n7359), .Y(N34934) );
  AND2X2 U15789 ( .A(N34933), .B(n8403), .Y(N34950) );
  MX4X1 U15790 ( .A(n7263), .B(n7261), .C(n7262), .D(n7260), .S0(n7357), .S1(
        n7359), .Y(N34933) );
  AND2X2 U15791 ( .A(N34932), .B(n8403), .Y(N34951) );
  MX4X1 U15792 ( .A(n7267), .B(n7265), .C(n7266), .D(n7264), .S0(n7357), .S1(
        n7359), .Y(N34932) );
  AND2X2 U15793 ( .A(N34931), .B(n8403), .Y(N34952) );
  MX4X1 U15794 ( .A(n7271), .B(n7269), .C(n7270), .D(n7268), .S0(n7357), .S1(
        n7359), .Y(N34931) );
  AND2X2 U15795 ( .A(N34930), .B(n8403), .Y(N34953) );
  MX4X1 U15796 ( .A(n7275), .B(n7273), .C(n7274), .D(n7272), .S0(n7357), .S1(
        n7359), .Y(N34930) );
  AND2X2 U15797 ( .A(N34929), .B(n8403), .Y(N34954) );
  MX4X1 U15798 ( .A(n7279), .B(n7277), .C(n7278), .D(n7276), .S0(n7357), .S1(
        n7359), .Y(N34929) );
  AND2X2 U15799 ( .A(N34928), .B(n8403), .Y(N34955) );
  MX4X1 U15800 ( .A(n7283), .B(n7281), .C(n7282), .D(n7280), .S0(n7357), .S1(
        n7359), .Y(N34928) );
  AND2X2 U15801 ( .A(N34927), .B(n8403), .Y(N34956) );
  MX4X1 U15802 ( .A(n7287), .B(n7285), .C(n7286), .D(n7284), .S0(n7357), .S1(
        n7359), .Y(N34927) );
  AND2X2 U15803 ( .A(N34926), .B(n8403), .Y(N34957) );
  MX4X1 U15804 ( .A(n7291), .B(n7289), .C(n7290), .D(n7288), .S0(n7357), .S1(
        n7359), .Y(N34926) );
  AND2X2 U15805 ( .A(N34925), .B(n8403), .Y(N34958) );
  MX4X1 U15806 ( .A(n7295), .B(n7293), .C(n7294), .D(n7292), .S0(n7357), .S1(
        n7359), .Y(N34925) );
  AND2X2 U15807 ( .A(N34924), .B(n8403), .Y(N34959) );
  MX4X1 U15808 ( .A(n7299), .B(n7297), .C(n7298), .D(n7296), .S0(n7357), .S1(
        n7359), .Y(N34924) );
  AND2X2 U15809 ( .A(N34923), .B(n8403), .Y(N34960) );
  MX4X1 U15810 ( .A(n7303), .B(n7301), .C(n7302), .D(n7300), .S0(n7357), .S1(
        n7359), .Y(N34923) );
  AND2X2 U15811 ( .A(N34922), .B(n8403), .Y(N34961) );
  MX4X1 U15812 ( .A(n7307), .B(n7305), .C(n7306), .D(n7304), .S0(n7358), .S1(
        n7360), .Y(N34922) );
  AND2X2 U15813 ( .A(N34921), .B(n8402), .Y(N34962) );
  MX4X1 U15814 ( .A(n7311), .B(n7309), .C(n7310), .D(n7308), .S0(n7358), .S1(
        n7360), .Y(N34921) );
  AND2X2 U15815 ( .A(N34920), .B(n8402), .Y(N34963) );
  MX4X1 U15816 ( .A(n7315), .B(n7313), .C(n7314), .D(n7312), .S0(n7358), .S1(
        n7360), .Y(N34920) );
  AND2X2 U15817 ( .A(N34919), .B(n8402), .Y(N34964) );
  MX4X1 U15818 ( .A(n7319), .B(n7317), .C(n7318), .D(n7316), .S0(n7358), .S1(
        n7360), .Y(N34919) );
  AND2X2 U15819 ( .A(N34918), .B(n8402), .Y(N34965) );
  MX4X1 U15820 ( .A(n7323), .B(n7321), .C(n7322), .D(n7320), .S0(n7358), .S1(
        n7360), .Y(N34918) );
  AND2X2 U15821 ( .A(N34917), .B(n8402), .Y(N34966) );
  MX4X1 U15822 ( .A(n7327), .B(n7325), .C(n7326), .D(n7324), .S0(n7358), .S1(
        n7360), .Y(N34917) );
  AND2X2 U15823 ( .A(N34916), .B(n8402), .Y(N34967) );
  MX4X1 U15824 ( .A(n7331), .B(n7329), .C(n7330), .D(n7328), .S0(n7358), .S1(
        n7360), .Y(N34916) );
  AND2X2 U15825 ( .A(N34915), .B(n8402), .Y(N34968) );
  MX4X1 U15826 ( .A(n7335), .B(n7333), .C(n7334), .D(n7332), .S0(n7358), .S1(
        n7360), .Y(N34915) );
  AND2X2 U15827 ( .A(N34914), .B(n8402), .Y(N34969) );
  MX4X1 U15828 ( .A(n7339), .B(n7337), .C(n7338), .D(n7336), .S0(n7358), .S1(
        n7360), .Y(N34914) );
  AND2X2 U15829 ( .A(N34913), .B(n8402), .Y(N34970) );
  MX4X1 U15830 ( .A(n7343), .B(n7341), .C(n7342), .D(n7340), .S0(n7358), .S1(
        n7360), .Y(N34913) );
  AND2X2 U15831 ( .A(N34912), .B(n8402), .Y(N34971) );
  MX4X1 U15832 ( .A(n7347), .B(n7345), .C(n7346), .D(n7344), .S0(
        outCount_next[3]), .S1(n7360), .Y(N34912) );
  AND2X2 U15833 ( .A(N34911), .B(n8402), .Y(N34972) );
  MX4X1 U15834 ( .A(n7351), .B(n7349), .C(n7350), .D(n7348), .S0(n7358), .S1(
        n7360), .Y(N34911) );
  AND2X2 U15835 ( .A(N34910), .B(n8402), .Y(N34973) );
  MX4X1 U15836 ( .A(n7355), .B(n7353), .C(n7354), .D(n7352), .S0(n7358), .S1(
        n7360), .Y(N34910) );
  NOR2X1 U15837 ( .A(n6995), .B(n5703), .Y(n2937) );
  NOR2X1 U15838 ( .A(n7004), .B(n5702), .Y(n2730) );
  NOR4X1 U15839 ( .A(n4900), .B(n4901), .C(n73), .D(n8404), .Y(n4894) );
  NAND2X1 U15840 ( .A(n76), .B(n75), .Y(n4901) );
  NAND4X1 U15841 ( .A(n80), .B(n79), .C(n78), .D(n77), .Y(n4900) );
  NAND2X1 U15842 ( .A(state[1]), .B(n6624), .Y(n161) );
  NAND4X1 U15843 ( .A(n4892), .B(n4893), .C(n4894), .D(n4895), .Y(n4883) );
  AND4X1 U15844 ( .A(n85), .B(n86), .C(n87), .D(n88), .Y(n4892) );
  AND4X1 U15845 ( .A(n81), .B(n82), .C(n83), .D(n84), .Y(n4893) );
  NOR4X1 U15846 ( .A(n4896), .B(n4897), .C(n4898), .D(n4899), .Y(n4895) );
  OAI22XL U15847 ( .A0(n4934), .A1(n7699), .B0(n8845), .B1(n216), .Y(n5739) );
  OAI22XL U15848 ( .A0(n4935), .A1(n7699), .B0(n8844), .B1(n216), .Y(n5740) );
  OAI22XL U15849 ( .A0(n4936), .A1(n7699), .B0(n8843), .B1(n216), .Y(n5741) );
  OAI22XL U15850 ( .A0(n4937), .A1(n7699), .B0(n8842), .B1(n216), .Y(n5742) );
  OAI22XL U15851 ( .A0(n4938), .A1(n7699), .B0(n8841), .B1(n216), .Y(n5743) );
  OAI22XL U15852 ( .A0(n4939), .A1(n7699), .B0(n8840), .B1(n216), .Y(n5744) );
  OAI22XL U15853 ( .A0(n4940), .A1(n7699), .B0(n8839), .B1(n216), .Y(n5745) );
  OAI22XL U15854 ( .A0(n4941), .A1(n7699), .B0(n8838), .B1(n216), .Y(n5746) );
  OAI22XL U15855 ( .A0(n4942), .A1(n7699), .B0(n8837), .B1(n216), .Y(n5747) );
  OAI22XL U15856 ( .A0(n4943), .A1(n7699), .B0(n8836), .B1(n216), .Y(n5748) );
  OAI22XL U15857 ( .A0(n4944), .A1(n7699), .B0(n8835), .B1(n216), .Y(n5749) );
  OAI22XL U15858 ( .A0(n4945), .A1(n6719), .B0(n8834), .B1(n216), .Y(n5750) );
  OAI22XL U15859 ( .A0(n4946), .A1(n6719), .B0(n8833), .B1(n216), .Y(n5751) );
  OAI22XL U15860 ( .A0(n4947), .A1(n6719), .B0(n8832), .B1(n216), .Y(n5752) );
  OAI22XL U15861 ( .A0(n4948), .A1(n6719), .B0(n8831), .B1(n216), .Y(n5753) );
  OAI22XL U15862 ( .A0(n4982), .A1(n7687), .B0(n8845), .B1(n219), .Y(n5787) );
  OAI22XL U15863 ( .A0(n4983), .A1(n7687), .B0(n8844), .B1(n219), .Y(n5788) );
  OAI22XL U15864 ( .A0(n4984), .A1(n7687), .B0(n8843), .B1(n219), .Y(n5789) );
  OAI22XL U15865 ( .A0(n4985), .A1(n7687), .B0(n8842), .B1(n219), .Y(n5790) );
  OAI22XL U15866 ( .A0(n4986), .A1(n7687), .B0(n8841), .B1(n219), .Y(n5791) );
  OAI22XL U15867 ( .A0(n4987), .A1(n7687), .B0(n8840), .B1(n219), .Y(n5792) );
  OAI22XL U15868 ( .A0(n4988), .A1(n7687), .B0(n8839), .B1(n219), .Y(n5793) );
  OAI22XL U15869 ( .A0(n4989), .A1(n7687), .B0(n8838), .B1(n219), .Y(n5794) );
  OAI22XL U15870 ( .A0(n4990), .A1(n7687), .B0(n8837), .B1(n219), .Y(n5795) );
  OAI22XL U15871 ( .A0(n4991), .A1(n7687), .B0(n8836), .B1(n219), .Y(n5796) );
  OAI22XL U15872 ( .A0(n4992), .A1(n7687), .B0(n8835), .B1(n219), .Y(n5797) );
  OAI22XL U15873 ( .A0(n4993), .A1(n7687), .B0(n8834), .B1(n219), .Y(n5798) );
  OAI22XL U15874 ( .A0(n4994), .A1(n7687), .B0(n8833), .B1(n219), .Y(n5799) );
  OAI22XL U15875 ( .A0(n4995), .A1(n7687), .B0(n8832), .B1(n219), .Y(n5800) );
  OAI22XL U15876 ( .A0(n4996), .A1(n6720), .B0(n8831), .B1(n219), .Y(n5801) );
  OAI22XL U15877 ( .A0(n5030), .A1(n7689), .B0(n8845), .B1(n223), .Y(n5835) );
  OAI22XL U15878 ( .A0(n5031), .A1(n7689), .B0(n8844), .B1(n223), .Y(n5836) );
  OAI22XL U15879 ( .A0(n5032), .A1(n7689), .B0(n8843), .B1(n223), .Y(n5837) );
  OAI22XL U15880 ( .A0(n5033), .A1(n7689), .B0(n8842), .B1(n223), .Y(n5838) );
  OAI22XL U15881 ( .A0(n5034), .A1(n7689), .B0(n8841), .B1(n223), .Y(n5839) );
  OAI22XL U15882 ( .A0(n5035), .A1(n7689), .B0(n8840), .B1(n223), .Y(n5840) );
  OAI22XL U15883 ( .A0(n5036), .A1(n7689), .B0(n8839), .B1(n223), .Y(n5841) );
  OAI22XL U15884 ( .A0(n5037), .A1(n7689), .B0(n8838), .B1(n223), .Y(n5842) );
  OAI22XL U15885 ( .A0(n5038), .A1(n7689), .B0(n8837), .B1(n223), .Y(n5843) );
  OAI22XL U15886 ( .A0(n5039), .A1(n7689), .B0(n8836), .B1(n223), .Y(n5844) );
  OAI22XL U15887 ( .A0(n5040), .A1(n7689), .B0(n8835), .B1(n223), .Y(n5845) );
  OAI22XL U15888 ( .A0(n5041), .A1(n6721), .B0(n8834), .B1(n223), .Y(n5846) );
  OAI22XL U15889 ( .A0(n5042), .A1(n6721), .B0(n8833), .B1(n223), .Y(n5847) );
  OAI22XL U15890 ( .A0(n5043), .A1(n6721), .B0(n8832), .B1(n223), .Y(n5848) );
  OAI22XL U15891 ( .A0(n5044), .A1(n6721), .B0(n8831), .B1(n223), .Y(n5849) );
  OAI22XL U15892 ( .A0(n5078), .A1(n7691), .B0(n8845), .B1(n227), .Y(n5883) );
  OAI22XL U15893 ( .A0(n5079), .A1(n7691), .B0(n8844), .B1(n227), .Y(n5884) );
  OAI22XL U15894 ( .A0(n5080), .A1(n7691), .B0(n8843), .B1(n227), .Y(n5885) );
  OAI22XL U15895 ( .A0(n5081), .A1(n7691), .B0(n8842), .B1(n227), .Y(n5886) );
  OAI22XL U15896 ( .A0(n5082), .A1(n7691), .B0(n8841), .B1(n227), .Y(n5887) );
  OAI22XL U15897 ( .A0(n5083), .A1(n7691), .B0(n8840), .B1(n227), .Y(n5888) );
  OAI22XL U15898 ( .A0(n5084), .A1(n7691), .B0(n8839), .B1(n227), .Y(n5889) );
  OAI22XL U15899 ( .A0(n5085), .A1(n7691), .B0(n8838), .B1(n227), .Y(n5890) );
  OAI22XL U15900 ( .A0(n5086), .A1(n7691), .B0(n8837), .B1(n227), .Y(n5891) );
  OAI22XL U15901 ( .A0(n5087), .A1(n7691), .B0(n8836), .B1(n227), .Y(n5892) );
  OAI22XL U15902 ( .A0(n5088), .A1(n7691), .B0(n8835), .B1(n227), .Y(n5893) );
  OAI22XL U15903 ( .A0(n5089), .A1(n7691), .B0(n8834), .B1(n227), .Y(n5894) );
  OAI22XL U15904 ( .A0(n5090), .A1(n7691), .B0(n8833), .B1(n227), .Y(n5895) );
  OAI22XL U15905 ( .A0(n5091), .A1(n7691), .B0(n8832), .B1(n227), .Y(n5896) );
  OAI22XL U15906 ( .A0(n5092), .A1(n6722), .B0(n8831), .B1(n227), .Y(n5897) );
  OAI22XL U15907 ( .A0(n5126), .A1(n7693), .B0(n8845), .B1(n231), .Y(n5931) );
  OAI22XL U15908 ( .A0(n5127), .A1(n7693), .B0(n8844), .B1(n231), .Y(n5932) );
  OAI22XL U15909 ( .A0(n5128), .A1(n7693), .B0(n8843), .B1(n231), .Y(n5933) );
  OAI22XL U15910 ( .A0(n5129), .A1(n7693), .B0(n8842), .B1(n231), .Y(n5934) );
  OAI22XL U15911 ( .A0(n5130), .A1(n7693), .B0(n8841), .B1(n231), .Y(n5935) );
  OAI22XL U15912 ( .A0(n5131), .A1(n7693), .B0(n8840), .B1(n231), .Y(n5936) );
  OAI22XL U15913 ( .A0(n5132), .A1(n7693), .B0(n8839), .B1(n231), .Y(n5937) );
  OAI22XL U15914 ( .A0(n5133), .A1(n7693), .B0(n8838), .B1(n231), .Y(n5938) );
  OAI22XL U15915 ( .A0(n5134), .A1(n7693), .B0(n8837), .B1(n231), .Y(n5939) );
  OAI22XL U15916 ( .A0(n5135), .A1(n7693), .B0(n8836), .B1(n231), .Y(n5940) );
  OAI22XL U15917 ( .A0(n5136), .A1(n7693), .B0(n8835), .B1(n231), .Y(n5941) );
  OAI22XL U15918 ( .A0(n5137), .A1(n6723), .B0(n8834), .B1(n231), .Y(n5942) );
  OAI22XL U15919 ( .A0(n5138), .A1(n6723), .B0(n8833), .B1(n231), .Y(n5943) );
  OAI22XL U15920 ( .A0(n5139), .A1(n6723), .B0(n8832), .B1(n231), .Y(n5944) );
  OAI22XL U15921 ( .A0(n5140), .A1(n6723), .B0(n8831), .B1(n231), .Y(n5945) );
  OAI22XL U15922 ( .A0(n5174), .A1(n7695), .B0(n8845), .B1(n235), .Y(n5979) );
  OAI22XL U15923 ( .A0(n5175), .A1(n7695), .B0(n8844), .B1(n235), .Y(n5980) );
  OAI22XL U15924 ( .A0(n5176), .A1(n7695), .B0(n8843), .B1(n235), .Y(n5981) );
  OAI22XL U15925 ( .A0(n5177), .A1(n7695), .B0(n8842), .B1(n235), .Y(n5982) );
  OAI22XL U15926 ( .A0(n5178), .A1(n7695), .B0(n8841), .B1(n235), .Y(n5983) );
  OAI22XL U15927 ( .A0(n5179), .A1(n7695), .B0(n8840), .B1(n235), .Y(n5984) );
  OAI22XL U15928 ( .A0(n5180), .A1(n7695), .B0(n8839), .B1(n235), .Y(n5985) );
  OAI22XL U15929 ( .A0(n5181), .A1(n7695), .B0(n8838), .B1(n235), .Y(n5986) );
  OAI22XL U15930 ( .A0(n5182), .A1(n7695), .B0(n8837), .B1(n235), .Y(n5987) );
  OAI22XL U15931 ( .A0(n5183), .A1(n7695), .B0(n8836), .B1(n235), .Y(n5988) );
  OAI22XL U15932 ( .A0(n5184), .A1(n7695), .B0(n8835), .B1(n235), .Y(n5989) );
  OAI22XL U15933 ( .A0(n5185), .A1(n6724), .B0(n8834), .B1(n235), .Y(n5990) );
  OAI22XL U15934 ( .A0(n5186), .A1(n6724), .B0(n8833), .B1(n235), .Y(n5991) );
  OAI22XL U15935 ( .A0(n5187), .A1(n6724), .B0(n8832), .B1(n235), .Y(n5992) );
  OAI22XL U15936 ( .A0(n5188), .A1(n6724), .B0(n8831), .B1(n235), .Y(n5993) );
  OAI22XL U15937 ( .A0(n5270), .A1(n7671), .B0(n8845), .B1(n184), .Y(n6075) );
  OAI22XL U15938 ( .A0(n5271), .A1(n7671), .B0(n8844), .B1(n184), .Y(n6076) );
  OAI22XL U15939 ( .A0(n5272), .A1(n7671), .B0(n8843), .B1(n184), .Y(n6077) );
  OAI22XL U15940 ( .A0(n5273), .A1(n7671), .B0(n8842), .B1(n184), .Y(n6078) );
  OAI22XL U15941 ( .A0(n5274), .A1(n7671), .B0(n8841), .B1(n184), .Y(n6079) );
  OAI22XL U15942 ( .A0(n5275), .A1(n7671), .B0(n8840), .B1(n184), .Y(n6080) );
  OAI22XL U15943 ( .A0(n5276), .A1(n7671), .B0(n8839), .B1(n184), .Y(n6081) );
  OAI22XL U15944 ( .A0(n5277), .A1(n7671), .B0(n8838), .B1(n184), .Y(n6082) );
  OAI22XL U15945 ( .A0(n5278), .A1(n7671), .B0(n8837), .B1(n184), .Y(n6083) );
  OAI22XL U15946 ( .A0(n5279), .A1(n7671), .B0(n8836), .B1(n184), .Y(n6084) );
  OAI22XL U15947 ( .A0(n5280), .A1(n7671), .B0(n8835), .B1(n184), .Y(n6085) );
  OAI22XL U15948 ( .A0(n5281), .A1(n6725), .B0(n8834), .B1(n184), .Y(n6086) );
  OAI22XL U15949 ( .A0(n5282), .A1(n6725), .B0(n8833), .B1(n184), .Y(n6087) );
  OAI22XL U15950 ( .A0(n5283), .A1(n6725), .B0(n8832), .B1(n184), .Y(n6088) );
  OAI22XL U15951 ( .A0(n5284), .A1(n6725), .B0(n8831), .B1(n184), .Y(n6089) );
  OAI22XL U15952 ( .A0(n5318), .A1(n7673), .B0(n8845), .B1(n188), .Y(n6123) );
  OAI22XL U15953 ( .A0(n5319), .A1(n7673), .B0(n8844), .B1(n188), .Y(n6124) );
  OAI22XL U15954 ( .A0(n5320), .A1(n7673), .B0(n8843), .B1(n188), .Y(n6125) );
  OAI22XL U15955 ( .A0(n5321), .A1(n7673), .B0(n8842), .B1(n188), .Y(n6126) );
  OAI22XL U15956 ( .A0(n5322), .A1(n7673), .B0(n8841), .B1(n188), .Y(n6127) );
  OAI22XL U15957 ( .A0(n5323), .A1(n7673), .B0(n8840), .B1(n188), .Y(n6128) );
  OAI22XL U15958 ( .A0(n5324), .A1(n7673), .B0(n8839), .B1(n188), .Y(n6129) );
  OAI22XL U15959 ( .A0(n5325), .A1(n7673), .B0(n8838), .B1(n188), .Y(n6130) );
  OAI22XL U15960 ( .A0(n5326), .A1(n7673), .B0(n8837), .B1(n188), .Y(n6131) );
  OAI22XL U15961 ( .A0(n5327), .A1(n7673), .B0(n8836), .B1(n188), .Y(n6132) );
  OAI22XL U15962 ( .A0(n5328), .A1(n7673), .B0(n8835), .B1(n188), .Y(n6133) );
  OAI22XL U15963 ( .A0(n5329), .A1(n6726), .B0(n8834), .B1(n188), .Y(n6134) );
  OAI22XL U15964 ( .A0(n5330), .A1(n6726), .B0(n8833), .B1(n188), .Y(n6135) );
  OAI22XL U15965 ( .A0(n5331), .A1(n6726), .B0(n8832), .B1(n188), .Y(n6136) );
  OAI22XL U15966 ( .A0(n5332), .A1(n6726), .B0(n8831), .B1(n188), .Y(n6137) );
  OAI22XL U15967 ( .A0(n5366), .A1(n7675), .B0(n8845), .B1(n192), .Y(n6171) );
  OAI22XL U15968 ( .A0(n5367), .A1(n7675), .B0(n8844), .B1(n192), .Y(n6172) );
  OAI22XL U15969 ( .A0(n5368), .A1(n7675), .B0(n8843), .B1(n192), .Y(n6173) );
  OAI22XL U15970 ( .A0(n5369), .A1(n7675), .B0(n8842), .B1(n192), .Y(n6174) );
  OAI22XL U15971 ( .A0(n5370), .A1(n7675), .B0(n8841), .B1(n192), .Y(n6175) );
  OAI22XL U15972 ( .A0(n5371), .A1(n7675), .B0(n8840), .B1(n192), .Y(n6176) );
  OAI22XL U15973 ( .A0(n5372), .A1(n7675), .B0(n8839), .B1(n192), .Y(n6177) );
  OAI22XL U15974 ( .A0(n5373), .A1(n7675), .B0(n8838), .B1(n192), .Y(n6178) );
  OAI22XL U15975 ( .A0(n5374), .A1(n7675), .B0(n8837), .B1(n192), .Y(n6179) );
  OAI22XL U15976 ( .A0(n5375), .A1(n7675), .B0(n8836), .B1(n192), .Y(n6180) );
  OAI22XL U15977 ( .A0(n5376), .A1(n7675), .B0(n8835), .B1(n192), .Y(n6181) );
  OAI22XL U15978 ( .A0(n5377), .A1(n7675), .B0(n8834), .B1(n192), .Y(n6182) );
  OAI22XL U15979 ( .A0(n5378), .A1(n7675), .B0(n8833), .B1(n192), .Y(n6183) );
  OAI22XL U15980 ( .A0(n5379), .A1(n7675), .B0(n8832), .B1(n192), .Y(n6184) );
  OAI22XL U15981 ( .A0(n5380), .A1(n6727), .B0(n8831), .B1(n192), .Y(n6185) );
  OAI22XL U15982 ( .A0(n5414), .A1(n7677), .B0(n8845), .B1(n196), .Y(n6219) );
  OAI22XL U15983 ( .A0(n5415), .A1(n7677), .B0(n8844), .B1(n196), .Y(n6220) );
  OAI22XL U15984 ( .A0(n5416), .A1(n7677), .B0(n8843), .B1(n196), .Y(n6221) );
  OAI22XL U15985 ( .A0(n5417), .A1(n7677), .B0(n8842), .B1(n196), .Y(n6222) );
  OAI22XL U15986 ( .A0(n5418), .A1(n7677), .B0(n8841), .B1(n196), .Y(n6223) );
  OAI22XL U15987 ( .A0(n5419), .A1(n7677), .B0(n8840), .B1(n196), .Y(n6224) );
  OAI22XL U15988 ( .A0(n5420), .A1(n7677), .B0(n8839), .B1(n196), .Y(n6225) );
  OAI22XL U15989 ( .A0(n5421), .A1(n7677), .B0(n8838), .B1(n196), .Y(n6226) );
  OAI22XL U15990 ( .A0(n5422), .A1(n7677), .B0(n8837), .B1(n196), .Y(n6227) );
  OAI22XL U15991 ( .A0(n5423), .A1(n7677), .B0(n8836), .B1(n196), .Y(n6228) );
  OAI22XL U15992 ( .A0(n5424), .A1(n7677), .B0(n8835), .B1(n196), .Y(n6229) );
  OAI22XL U15993 ( .A0(n5425), .A1(n6728), .B0(n8834), .B1(n196), .Y(n6230) );
  OAI22XL U15994 ( .A0(n5426), .A1(n6728), .B0(n8833), .B1(n196), .Y(n6231) );
  OAI22XL U15995 ( .A0(n5427), .A1(n6728), .B0(n8832), .B1(n196), .Y(n6232) );
  OAI22XL U15996 ( .A0(n5428), .A1(n6728), .B0(n8831), .B1(n196), .Y(n6233) );
  OAI22XL U15997 ( .A0(n5462), .A1(n7679), .B0(n8845), .B1(n200), .Y(n6267) );
  OAI22XL U15998 ( .A0(n5463), .A1(n7679), .B0(n8844), .B1(n200), .Y(n6268) );
  OAI22XL U15999 ( .A0(n5464), .A1(n7679), .B0(n8843), .B1(n200), .Y(n6269) );
  OAI22XL U16000 ( .A0(n5465), .A1(n7679), .B0(n8842), .B1(n200), .Y(n6270) );
  OAI22XL U16001 ( .A0(n5466), .A1(n7679), .B0(n8841), .B1(n200), .Y(n6271) );
  OAI22XL U16002 ( .A0(n5467), .A1(n7679), .B0(n8840), .B1(n200), .Y(n6272) );
  OAI22XL U16003 ( .A0(n5468), .A1(n7679), .B0(n8839), .B1(n200), .Y(n6273) );
  OAI22XL U16004 ( .A0(n5469), .A1(n7679), .B0(n8838), .B1(n200), .Y(n6274) );
  OAI22XL U16005 ( .A0(n5470), .A1(n7679), .B0(n8837), .B1(n200), .Y(n6275) );
  OAI22XL U16006 ( .A0(n5471), .A1(n7679), .B0(n8836), .B1(n200), .Y(n6276) );
  OAI22XL U16007 ( .A0(n5472), .A1(n7679), .B0(n8835), .B1(n200), .Y(n6277) );
  OAI22XL U16008 ( .A0(n5473), .A1(n7679), .B0(n8834), .B1(n200), .Y(n6278) );
  OAI22XL U16009 ( .A0(n5474), .A1(n7679), .B0(n8833), .B1(n200), .Y(n6279) );
  OAI22XL U16010 ( .A0(n5475), .A1(n7679), .B0(n8832), .B1(n200), .Y(n6280) );
  OAI22XL U16011 ( .A0(n5476), .A1(n6729), .B0(n8831), .B1(n200), .Y(n6281) );
  OAI22XL U16012 ( .A0(n5510), .A1(n7681), .B0(n8845), .B1(n204), .Y(n6315) );
  OAI22XL U16013 ( .A0(n5511), .A1(n7681), .B0(n8844), .B1(n204), .Y(n6316) );
  OAI22XL U16014 ( .A0(n5512), .A1(n7681), .B0(n8843), .B1(n204), .Y(n6317) );
  OAI22XL U16015 ( .A0(n5513), .A1(n7681), .B0(n8842), .B1(n204), .Y(n6318) );
  OAI22XL U16016 ( .A0(n5514), .A1(n7681), .B0(n8841), .B1(n204), .Y(n6319) );
  OAI22XL U16017 ( .A0(n5515), .A1(n7681), .B0(n8840), .B1(n204), .Y(n6320) );
  OAI22XL U16018 ( .A0(n5516), .A1(n7681), .B0(n8839), .B1(n204), .Y(n6321) );
  OAI22XL U16019 ( .A0(n5517), .A1(n7681), .B0(n8838), .B1(n204), .Y(n6322) );
  OAI22XL U16020 ( .A0(n5518), .A1(n7681), .B0(n8837), .B1(n204), .Y(n6323) );
  OAI22XL U16021 ( .A0(n5519), .A1(n7681), .B0(n8836), .B1(n204), .Y(n6324) );
  OAI22XL U16022 ( .A0(n5520), .A1(n7681), .B0(n8835), .B1(n204), .Y(n6325) );
  OAI22XL U16023 ( .A0(n5521), .A1(n6730), .B0(n8834), .B1(n204), .Y(n6326) );
  OAI22XL U16024 ( .A0(n5522), .A1(n6730), .B0(n8833), .B1(n204), .Y(n6327) );
  OAI22XL U16025 ( .A0(n5523), .A1(n6730), .B0(n8832), .B1(n204), .Y(n6328) );
  OAI22XL U16026 ( .A0(n5524), .A1(n6730), .B0(n8831), .B1(n204), .Y(n6329) );
  OAI22XL U16027 ( .A0(n5558), .A1(n7683), .B0(n8845), .B1(n208), .Y(n6363) );
  OAI22XL U16028 ( .A0(n5559), .A1(n7683), .B0(n8844), .B1(n208), .Y(n6364) );
  OAI22XL U16029 ( .A0(n5560), .A1(n7683), .B0(n8843), .B1(n208), .Y(n6365) );
  OAI22XL U16030 ( .A0(n5561), .A1(n7683), .B0(n8842), .B1(n208), .Y(n6366) );
  OAI22XL U16031 ( .A0(n5562), .A1(n7683), .B0(n8841), .B1(n208), .Y(n6367) );
  OAI22XL U16032 ( .A0(n5563), .A1(n7683), .B0(n8840), .B1(n208), .Y(n6368) );
  OAI22XL U16033 ( .A0(n5564), .A1(n7683), .B0(n8839), .B1(n208), .Y(n6369) );
  OAI22XL U16034 ( .A0(n5565), .A1(n7683), .B0(n8838), .B1(n208), .Y(n6370) );
  OAI22XL U16035 ( .A0(n5566), .A1(n7683), .B0(n8837), .B1(n208), .Y(n6371) );
  OAI22XL U16036 ( .A0(n5567), .A1(n7683), .B0(n8836), .B1(n208), .Y(n6372) );
  OAI22XL U16037 ( .A0(n5568), .A1(n7683), .B0(n8835), .B1(n208), .Y(n6373) );
  OAI22XL U16038 ( .A0(n5569), .A1(n6731), .B0(n8834), .B1(n208), .Y(n6374) );
  OAI22XL U16039 ( .A0(n5570), .A1(n6731), .B0(n8833), .B1(n208), .Y(n6375) );
  OAI22XL U16040 ( .A0(n5571), .A1(n6731), .B0(n8832), .B1(n208), .Y(n6376) );
  OAI22XL U16041 ( .A0(n5572), .A1(n6731), .B0(n8831), .B1(n208), .Y(n6377) );
  OAI22XL U16042 ( .A0(n5606), .A1(n7685), .B0(n8845), .B1(n212), .Y(n6411) );
  OAI22XL U16043 ( .A0(n5607), .A1(n7685), .B0(n8844), .B1(n212), .Y(n6412) );
  OAI22XL U16044 ( .A0(n5608), .A1(n7685), .B0(n8843), .B1(n212), .Y(n6413) );
  OAI22XL U16045 ( .A0(n5609), .A1(n7685), .B0(n8842), .B1(n212), .Y(n6414) );
  OAI22XL U16046 ( .A0(n5610), .A1(n7685), .B0(n8841), .B1(n212), .Y(n6415) );
  OAI22XL U16047 ( .A0(n5611), .A1(n7685), .B0(n8840), .B1(n212), .Y(n6416) );
  OAI22XL U16048 ( .A0(n5612), .A1(n7685), .B0(n8839), .B1(n212), .Y(n6417) );
  OAI22XL U16049 ( .A0(n5613), .A1(n7685), .B0(n8838), .B1(n212), .Y(n6418) );
  OAI22XL U16050 ( .A0(n5614), .A1(n7685), .B0(n8837), .B1(n212), .Y(n6419) );
  OAI22XL U16051 ( .A0(n5615), .A1(n7685), .B0(n8836), .B1(n212), .Y(n6420) );
  OAI22XL U16052 ( .A0(n5616), .A1(n7685), .B0(n8835), .B1(n212), .Y(n6421) );
  OAI22XL U16053 ( .A0(n5617), .A1(n6732), .B0(n8834), .B1(n212), .Y(n6422) );
  OAI22XL U16054 ( .A0(n5618), .A1(n6732), .B0(n8833), .B1(n212), .Y(n6423) );
  OAI22XL U16055 ( .A0(n5619), .A1(n6732), .B0(n8832), .B1(n212), .Y(n6424) );
  OAI22XL U16056 ( .A0(n5620), .A1(n6732), .B0(n8831), .B1(n212), .Y(n6425) );
  OAI22XL U16057 ( .A0(n5654), .A1(n7697), .B0(n8845), .B1(n239), .Y(n6459) );
  OAI22XL U16058 ( .A0(n5655), .A1(n7697), .B0(n8844), .B1(n239), .Y(n6460) );
  OAI22XL U16059 ( .A0(n5656), .A1(n7697), .B0(n8843), .B1(n239), .Y(n6461) );
  OAI22XL U16060 ( .A0(n5657), .A1(n7697), .B0(n8842), .B1(n239), .Y(n6462) );
  OAI22XL U16061 ( .A0(n5658), .A1(n7697), .B0(n8841), .B1(n239), .Y(n6463) );
  OAI22XL U16062 ( .A0(n5659), .A1(n7697), .B0(n8840), .B1(n239), .Y(n6464) );
  OAI22XL U16063 ( .A0(n5660), .A1(n7697), .B0(n8839), .B1(n239), .Y(n6465) );
  OAI22XL U16064 ( .A0(n5661), .A1(n7697), .B0(n8838), .B1(n239), .Y(n6466) );
  OAI22XL U16065 ( .A0(n5662), .A1(n7697), .B0(n8837), .B1(n239), .Y(n6467) );
  OAI22XL U16066 ( .A0(n5663), .A1(n7697), .B0(n8836), .B1(n239), .Y(n6468) );
  OAI22XL U16067 ( .A0(n5664), .A1(n7697), .B0(n8835), .B1(n239), .Y(n6469) );
  OAI22XL U16068 ( .A0(n5665), .A1(n6733), .B0(n8834), .B1(n239), .Y(n6470) );
  OAI22XL U16069 ( .A0(n5666), .A1(n6733), .B0(n8833), .B1(n239), .Y(n6471) );
  OAI22XL U16070 ( .A0(n5667), .A1(n6733), .B0(n8832), .B1(n239), .Y(n6472) );
  OAI22XL U16071 ( .A0(n5668), .A1(n6733), .B0(n8831), .B1(n239), .Y(n6473) );
  OAI22XL U16072 ( .A0(n5222), .A1(n7669), .B0(n165), .B1(n8845), .Y(n6027) );
  OAI22XL U16073 ( .A0(n5223), .A1(n7669), .B0(n165), .B1(n8844), .Y(n6028) );
  OAI22XL U16074 ( .A0(n5224), .A1(n7669), .B0(n165), .B1(n8843), .Y(n6029) );
  OAI22XL U16075 ( .A0(n5225), .A1(n7669), .B0(n165), .B1(n8842), .Y(n6030) );
  OAI22XL U16076 ( .A0(n5226), .A1(n7669), .B0(n165), .B1(n8841), .Y(n6031) );
  OAI22XL U16077 ( .A0(n5227), .A1(n7669), .B0(n165), .B1(n8840), .Y(n6032) );
  OAI22XL U16078 ( .A0(n5228), .A1(n7669), .B0(n165), .B1(n8839), .Y(n6033) );
  OAI22XL U16079 ( .A0(n5229), .A1(n7669), .B0(n165), .B1(n8838), .Y(n6034) );
  OAI22XL U16080 ( .A0(n5230), .A1(n7669), .B0(n165), .B1(n8837), .Y(n6035) );
  OAI22XL U16081 ( .A0(n5231), .A1(n7669), .B0(n165), .B1(n8836), .Y(n6036) );
  OAI22XL U16082 ( .A0(n5232), .A1(n7669), .B0(n165), .B1(n8835), .Y(n6037) );
  OAI22XL U16083 ( .A0(n5233), .A1(n6734), .B0(n165), .B1(n8834), .Y(n6038) );
  OAI22XL U16084 ( .A0(n5234), .A1(n6734), .B0(n165), .B1(n8833), .Y(n6039) );
  OAI22XL U16085 ( .A0(n5235), .A1(n6734), .B0(n165), .B1(n8832), .Y(n6040) );
  OAI22XL U16086 ( .A0(n5236), .A1(n6734), .B0(n165), .B1(n8831), .Y(n6041) );
  NAND4X1 U16087 ( .A(n6738), .B(n8853), .C(n4933), .D(n4932), .Y(n252) );
  NOR2X1 U16088 ( .A(n4929), .B(n4927), .Y(n6738) );
  CLKBUFX3 U16089 ( .A(N35189), .Y(n8405) );
  NAND4X1 U16090 ( .A(n74), .B(n5701), .C(n2524), .D(n101), .Y(n4899) );
  NAND4X1 U16091 ( .A(n100), .B(n99), .C(n98), .D(n97), .Y(n4898) );
  NAND4X1 U16092 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n4897) );
  NAND4X1 U16093 ( .A(n92), .B(n91), .C(n90), .D(n89), .Y(n4896) );
  AND4X1 U16094 ( .A(n4931), .B(n4930), .C(n4928), .D(n4926), .Y(n255) );
  AND4X1 U16095 ( .A(n4917), .B(n4916), .C(n4915), .D(n4914), .Y(n251) );
  AND4X1 U16096 ( .A(n4925), .B(n4924), .C(n4923), .D(n4922), .Y(n254) );
  AND4X1 U16097 ( .A(n4913), .B(n4912), .C(n4911), .D(n4910), .Y(n250) );
  AND4X1 U16098 ( .A(n4909), .B(n4908), .C(n4907), .D(n4906), .Y(n249) );
  AND4X1 U16099 ( .A(n4921), .B(n4920), .C(n4919), .D(n4918), .Y(n253) );
  AND4X1 U16100 ( .A(n4905), .B(n4904), .C(n4903), .D(n4902), .Y(n248) );
  CLKINVX1 U16101 ( .A(\xArray[4][42] ), .Y(n9057) );
  CLKINVX1 U16102 ( .A(\xArray[4][43] ), .Y(n9049) );
  CLKINVX1 U16103 ( .A(\xArray[4][44] ), .Y(n9041) );
  CLKINVX1 U16104 ( .A(\xArray[4][45] ), .Y(n9033) );
  CLKINVX1 U16105 ( .A(\xArray[4][46] ), .Y(n9025) );
  CLKINVX1 U16106 ( .A(\xArray[4][47] ), .Y(n9017) );
  CLKINVX1 U16107 ( .A(\xArray[4][48] ), .Y(n9009) );
  CLKINVX1 U16108 ( .A(\xArray[4][49] ), .Y(n9001) );
  CLKINVX1 U16109 ( .A(\xArray[4][50] ), .Y(n8993) );
  CLKINVX1 U16110 ( .A(\xArray[4][51] ), .Y(n8985) );
  CLKINVX1 U16111 ( .A(\xArray[4][52] ), .Y(n8977) );
  CLKINVX1 U16112 ( .A(\xArray[4][53] ), .Y(n8969) );
  CLKINVX1 U16113 ( .A(\xArray[4][54] ), .Y(n8961) );
  CLKINVX1 U16114 ( .A(\xArray[4][55] ), .Y(n8953) );
  CLKINVX1 U16115 ( .A(\xArray[4][56] ), .Y(n8945) );
  CLKINVX1 U16116 ( .A(\xArray[4][57] ), .Y(n8937) );
  CLKINVX1 U16117 ( .A(\xArray[4][58] ), .Y(n8929) );
  CLKINVX1 U16118 ( .A(\xArray[4][59] ), .Y(n8921) );
  CLKINVX1 U16119 ( .A(\xArray[4][60] ), .Y(n8913) );
  CLKINVX1 U16120 ( .A(\xArray[4][61] ), .Y(n8905) );
  CLKINVX1 U16121 ( .A(\xArray[4][62] ), .Y(n8897) );
  CLKINVX1 U16122 ( .A(\xArray[4][63] ), .Y(n8889) );
  CLKINVX1 U16123 ( .A(\xArray[15][42] ), .Y(n9055) );
  CLKINVX1 U16124 ( .A(\xArray[15][43] ), .Y(n9047) );
  CLKINVX1 U16125 ( .A(\xArray[15][44] ), .Y(n9039) );
  CLKINVX1 U16126 ( .A(\xArray[15][45] ), .Y(n9031) );
  CLKINVX1 U16127 ( .A(\xArray[15][46] ), .Y(n9023) );
  CLKINVX1 U16128 ( .A(\xArray[15][47] ), .Y(n9015) );
  CLKINVX1 U16129 ( .A(\xArray[15][48] ), .Y(n9007) );
  CLKINVX1 U16130 ( .A(\xArray[15][49] ), .Y(n8999) );
  CLKINVX1 U16131 ( .A(\xArray[15][50] ), .Y(n8991) );
  CLKINVX1 U16132 ( .A(\xArray[15][51] ), .Y(n8983) );
  CLKINVX1 U16133 ( .A(\xArray[15][52] ), .Y(n8975) );
  CLKINVX1 U16134 ( .A(\xArray[15][53] ), .Y(n8967) );
  CLKINVX1 U16135 ( .A(\xArray[15][54] ), .Y(n8959) );
  CLKINVX1 U16136 ( .A(\xArray[15][55] ), .Y(n8951) );
  CLKINVX1 U16137 ( .A(\xArray[15][56] ), .Y(n8943) );
  CLKINVX1 U16138 ( .A(\xArray[15][57] ), .Y(n8935) );
  CLKINVX1 U16139 ( .A(\xArray[15][58] ), .Y(n8927) );
  CLKINVX1 U16140 ( .A(\xArray[15][59] ), .Y(n8919) );
  CLKINVX1 U16141 ( .A(\xArray[15][60] ), .Y(n8911) );
  CLKINVX1 U16142 ( .A(\xArray[15][61] ), .Y(n8903) );
  CLKINVX1 U16143 ( .A(\xArray[15][62] ), .Y(n8895) );
  CLKINVX1 U16144 ( .A(\xArray[15][63] ), .Y(n8887) );
  MX4X2 U16145 ( .A(n7011), .B(n7009), .C(n7010), .D(n7008), .S0(n7224), .S1(
        n7223), .Y(N28880) );
  MX4X2 U16146 ( .A(n7175), .B(n7173), .C(n7174), .D(n7172), .S0(n7226), .S1(
        N1763), .Y(N28839) );
  MX4X2 U16147 ( .A(n7179), .B(n7177), .C(n7178), .D(n7176), .S0(n7226), .S1(
        N1763), .Y(N28838) );
  MX4X2 U16148 ( .A(n7183), .B(n7181), .C(n7182), .D(n7180), .S0(n7226), .S1(
        N1763), .Y(N28837) );
  MX4X2 U16149 ( .A(n7187), .B(n7185), .C(n7186), .D(n7184), .S0(n7226), .S1(
        N1763), .Y(N28836) );
  MX4X2 U16150 ( .A(n7191), .B(n7189), .C(n7190), .D(n7188), .S0(n8407), .S1(
        N1763), .Y(N28835) );
  MX4X2 U16151 ( .A(n7199), .B(n7197), .C(n7198), .D(n7196), .S0(n8407), .S1(
        N1763), .Y(N28833) );
  OAI221X4 U16152 ( .A0(n8309), .A1(n1292), .B0(n7716), .B1(n1548), .C0(n1549), 
        .Y(N33834) );
  OAI221X4 U16153 ( .A0(n8312), .A1(n1548), .B0(n7719), .B1(n1550), .C0(n1741), 
        .Y(N33770) );
  OAI211X4 U16154 ( .A0(n7751), .A1(n1548), .B0(n2315), .C0(n2316), .Y(N33706)
         );
  OAI221X4 U16155 ( .A0(n8317), .A1(n782), .B0(n7723), .B1(n780), .C0(n973), 
        .Y(N33962) );
  OAI221X4 U16156 ( .A0(n8312), .A1(n1287), .B0(n7716), .B1(n1544), .C0(n1545), 
        .Y(N33835) );
  NOR3X1 U16157 ( .A(iCount[21]), .B(iCount[23]), .C(iCount[22]), .Y(n8418) );
  NOR3X1 U16158 ( .A(iCount[24]), .B(iCount[26]), .C(iCount[25]), .Y(n8417) );
  NOR3X1 U16159 ( .A(iCount[27]), .B(iCount[29]), .C(iCount[28]), .Y(n8416) );
  NOR4X1 U16160 ( .A(iCount[9]), .B(iCount[8]), .C(iCount[31]), .D(iCount[30]), 
        .Y(n8415) );
  NAND4X1 U16161 ( .A(n8418), .B(n8417), .C(n8416), .D(n8415), .Y(n8425) );
  OR2X1 U16162 ( .A(iCount[5]), .B(iCount[4]), .Y(n8419) );
  AOI211X1 U16163 ( .A0(n8419), .A1(iCount[6]), .B0(iCount[7]), .C0(iCount[10]), .Y(n8423) );
  NOR3X1 U16164 ( .A(iCount[11]), .B(iCount[13]), .C(iCount[12]), .Y(n8422) );
  NOR3X1 U16165 ( .A(iCount[14]), .B(iCount[16]), .C(iCount[15]), .Y(n8421) );
  NOR4X1 U16166 ( .A(iCount[20]), .B(iCount[19]), .C(iCount[18]), .D(
        iCount[17]), .Y(n8420) );
  NAND4X1 U16167 ( .A(n8423), .B(n8422), .C(n8421), .D(n8420), .Y(n8424) );
  NOR3X1 U16168 ( .A(xCount[23]), .B(xCount[25]), .C(xCount[24]), .Y(n8429) );
  NOR4X1 U16169 ( .A(xCount[29]), .B(xCount[28]), .C(xCount[27]), .D(
        xCount[26]), .Y(n8428) );
  NOR4X1 U16170 ( .A(xCount[5]), .B(xCount[4]), .C(xCount[31]), .D(xCount[30]), 
        .Y(n8427) );
  NOR4X1 U16171 ( .A(xCount[9]), .B(xCount[8]), .C(xCount[7]), .D(xCount[6]), 
        .Y(n8426) );
  NAND4X1 U16172 ( .A(n8429), .B(n8428), .C(n8427), .D(n8426), .Y(n8436) );
  NOR3X1 U16173 ( .A(n8430), .B(xCount[11]), .C(xCount[10]), .Y(n8434) );
  NOR4X1 U16174 ( .A(xCount[15]), .B(xCount[14]), .C(xCount[13]), .D(
        xCount[12]), .Y(n8433) );
  NOR3X1 U16175 ( .A(xCount[16]), .B(xCount[18]), .C(xCount[17]), .Y(n8432) );
  NOR4X1 U16176 ( .A(xCount[22]), .B(xCount[21]), .C(xCount[20]), .D(
        xCount[19]), .Y(n8431) );
  NAND4X1 U16177 ( .A(n8434), .B(n8433), .C(n8432), .D(n8431), .Y(n8435) );
  NOR2X1 U16178 ( .A(n8436), .B(n8435), .Y(N34983) );
  NOR3X1 U16179 ( .A(outCount[23]), .B(outCount[25]), .C(outCount[24]), .Y(
        n8440) );
  NOR4X1 U16180 ( .A(outCount[29]), .B(outCount[28]), .C(outCount[27]), .D(
        outCount[26]), .Y(n8439) );
  NOR4X1 U16181 ( .A(outCount[5]), .B(outCount[4]), .C(outCount[31]), .D(
        outCount[30]), .Y(n8438) );
  NOR4X1 U16182 ( .A(outCount[9]), .B(outCount[8]), .C(outCount[7]), .D(
        outCount[6]), .Y(n8437) );
  NAND4X1 U16183 ( .A(n8440), .B(n8439), .C(n8438), .D(n8437), .Y(n8447) );
  AND4X1 U16184 ( .A(outCount[3]), .B(outCount[2]), .C(outCount[1]), .D(
        outCount[0]), .Y(n8441) );
  NOR3X1 U16185 ( .A(n8441), .B(outCount[11]), .C(outCount[10]), .Y(n8445) );
  NOR4X1 U16186 ( .A(outCount[15]), .B(outCount[14]), .C(outCount[13]), .D(
        outCount[12]), .Y(n8444) );
  NOR3X1 U16187 ( .A(outCount[16]), .B(outCount[18]), .C(outCount[17]), .Y(
        n8443) );
  NOR4X1 U16188 ( .A(outCount[22]), .B(outCount[21]), .C(outCount[20]), .D(
        outCount[19]), .Y(n8442) );
  NAND4X1 U16189 ( .A(n8445), .B(n8444), .C(n8443), .D(n8442), .Y(n8446) );
endmodule

